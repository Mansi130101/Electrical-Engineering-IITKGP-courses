CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
177209362 0
0
6 Title:
5 Name:
0
0
0
12
2 +V
167 440 108 0 1 3
0 21
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 74LS273
150 353 262 0 18 37
0 21 20 35 34 33 32 7 8 9
10 36 37 38 39 6 5 4 3
0
0 0 13024 270
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
4441 0 0
0
0
10 Ascii Key~
169 330 48 0 11 12
0 25 24 23 22 40 41 42 11 0
0 56
0
0 0 4640 512
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3618 0 0
0
0
6 74LS83
105 296 329 0 14 29
0 6 5 4 3 7 8 9 10 2
31 30 29 28 19
0
0 0 13024 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
9 CA 7-Seg~
184 150 410 0 18 19
10 12 13 14 15 17 16 18 43 27
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-62 -24 -27 -16
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
7 Buffer~
58 351 87 0 2 22
0 11 20
0
0 0 608 270
4 4050
-14 -19 14 -11
3 U3A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
7734 0 0
0
0
2 +V
167 150 321 0 1 3
0 26
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 74LS273
150 352 156 0 18 37
0 21 20 44 45 46 47 22 23 24
25 35 34 33 32 7 8 9 10
0
0 0 13024 270
7 74LS273
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
7 Ground~
168 253 291 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
14 Logic Display~
6 222 346 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
6 74LS47
187 266 414 0 14 29
0 31 30 29 28 48 49 18 16 17
15 14 13 12 50
0
0 0 13024 270
6 74LS47
-21 -60 21 -52
2 U1
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
9 Resistor~
219 150 347 0 4 5
0 27 26 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
40
18 4 3 0 0 0 0 2 4 0 0 2
307 299
307 299
17 3 4 0 0 0 0 2 4 0 0 2
316 299
316 299
16 2 5 0 0 0 0 2 4 0 0 2
325 299
325 299
15 1 6 0 0 0 0 2 4 0 0 2
334 299
334 299
5 0 7 0 0 8320 0 4 0 0 36 4
298 299
294 299
294 219
334 219
6 0 8 0 0 4224 0 4 0 0 35 3
289 299
289 210
325 210
7 0 9 0 0 4224 0 4 0 0 34 3
280 299
280 200
316 200
8 18 10 0 0 4224 0 4 8 0 0 3
271 299
271 193
306 193
1 8 11 0 0 0 0 6 3 0 0 2
351 72
351 72
13 1 12 0 0 8320 0 11 5 0 0 4
253 451
253 515
129 515
129 446
2 12 13 0 0 8320 0 5 11 0 0 4
135 446
135 505
262 505
262 451
3 11 14 0 0 8320 0 5 11 0 0 4
141 446
141 495
271 495
271 451
4 10 15 0 0 8320 0 5 11 0 0 4
147 446
147 485
280 485
280 451
6 8 16 0 0 8320 0 5 11 0 0 4
159 446
159 467
298 467
298 451
5 9 17 0 0 8320 0 5 11 0 0 4
153 446
153 476
289 476
289 451
7 7 18 0 0 8320 0 5 11 0 0 4
165 446
165 459
307 459
307 451
1 14 19 0 0 4224 0 10 4 0 0 3
222 364
253 364
253 363
2 0 20 0 0 12416 0 2 0 0 21 8
379 235
379 193
424 193
424 104
378 104
378 111
378 111
378 103
1 1 21 0 0 4224 0 1 2 0 0 3
440 117
440 229
388 229
1 1 21 0 0 0 0 8 1 0 0 4
387 123
387 119
440 119
440 117
2 2 20 0 0 0 0 8 6 0 0 4
378 129
378 103
351 103
351 102
4 7 22 0 0 4224 0 3 8 0 0 4
327 72
327 115
333 115
333 129
3 8 23 0 0 4224 0 3 8 0 0 4
321 72
321 115
324 115
324 129
2 9 24 0 0 4224 0 3 8 0 0 2
315 72
315 129
1 10 25 0 0 4224 0 3 8 0 0 4
309 72
309 115
306 115
306 129
1 2 26 0 0 12416 0 7 12 0 0 4
150 330
150 336
150 336
150 329
1 9 27 0 0 4224 0 12 5 0 0 4
150 365
150 376
150 376
150 374
1 9 2 0 0 4224 0 9 4 0 0 4
253 299
253 296
253 296
253 299
4 13 28 0 0 4224 0 11 4 0 0 4
280 381
280 355
280 355
280 363
3 12 29 0 0 4224 0 11 4 0 0 4
289 381
289 355
289 355
289 363
2 11 30 0 0 4224 0 11 4 0 0 4
298 381
298 355
298 355
298 363
1 10 31 0 0 4224 0 11 4 0 0 4
307 381
307 355
307 355
307 363
10 18 10 0 0 0 0 2 8 0 0 3
307 235
307 193
306 193
9 17 9 0 0 0 0 2 8 0 0 3
316 235
316 193
315 193
8 16 8 0 0 0 0 2 8 0 0 3
325 235
325 193
324 193
7 15 7 0 0 0 0 2 8 0 0 3
334 235
334 193
333 193
6 14 32 0 0 4224 0 2 8 0 0 3
343 235
343 193
342 193
5 13 33 0 0 4224 0 2 8 0 0 3
352 235
352 193
351 193
4 12 34 0 0 4224 0 2 8 0 0 3
361 235
361 193
360 193
3 11 35 0 0 4224 0 2 8 0 0 3
370 235
370 193
369 193
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 269
503 179 759 363
513 187 761 331
269 Here an one single digit adder 
is made. It outputs the sum of 
the last 2 subsequent digits 
entered as input to ASCII Key 
(used due to stroke providing 
input to the 8 bit register-
74LS273 ). Output is displayed 
with the help of 7 segment 
display.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
4.53041e-315 0 4.53041e-315 0 4.53041e-315 4.53041e-315
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
