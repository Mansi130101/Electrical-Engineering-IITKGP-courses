CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 80 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
177209362 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 233 211 0 1 11
0 3
0
0 0 21360 512
2 0V
2 -18 16 -10
2 V5
-9 9 5 17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 19 331 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
7 Buffer~
58 421 321 0 2 22
0 9 8
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U9B
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 4 0
1 U
3618 0 0
0
0
7 Buffer~
58 422 363 0 2 22
0 6 7
0
0 0 624 90
4 4050
-14 -19 14 -11
3 U9A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 4 0
1 U
6153 0 0
0
0
5 7415~
219 365 451 0 4 22
0 8 7 6 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
5394 0 0
0
0
9 Inverter~
13 418 415 0 2 22
0 10 6
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6A
-23 -7 -2 1
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
7734 0 0
0
0
7 Ground~
168 194 129 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
2 +V
167 64 234 0 1 3
0 17
0
0 0 54256 0
2 5V
-24 11 -10 19
2 V2
-22 0 -8 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
7 Ground~
168 64 380 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 145 291 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
6 1K RAM
79 192 321 0 20 41
0 2 2 2 2 2 2 26 25 24
23 36 37 38 39 11 12 13 14 2
15
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U5
-7 57 7 65
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
10 Ascii Key~
169 469 410 0 11 12
0 22 21 20 19 40 41 42 10 0
0 63
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
8903 0 0
0
0
7 74LS374
66 455 496 0 37 37
0 43 19 44 20 45 21 46 22 47
11 48 12 49 13 50 14 5 6 0
0 0 0 0 0 0 0 0 0 0
2 1 2 1 2 1 2 1
0
0 0 13040 782
7 74LS374
-24 -60 25 -52
2 U4
48 -4 62 4
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
7 74LS193
137 102 330 0 14 29
0 16 17 17 4 2 2 2 2 51
52 26 25 24 23
0
0 0 13040 0
7 74LS193
-24 -51 25 -43
2 U3
-7 -55 7 -47
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
7 74LS157
122 155 171 0 14 29
0 3 18 5 53 54 17 5 55 56
2 16 57 15 58
0
0 0 13040 180
7 74LS157
-24 -60 25 -52
2 U2
-13 -61 1 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Pulser~
4 69 98 0 10 12
0 59 60 18 61 0 0 5 5 3
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
9 CA 7-Seg~
184 68 640 0 18 19
10 29 30 31 32 34 33 35 62 28
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-62 -24 -27 -16
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
2 +V
167 68 560 0 1 3
0 27
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6671 0 0
0
0
6 74LS47
187 186 637 0 14 29
0 11 12 13 14 63 64 35 33 34
32 31 30 29 65
0
0 0 13040 782
6 74LS47
-21 -60 21 -52
2 U1
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
9 Resistor~
219 68 587 0 4 5
0 28 27 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
55
1 1 3 0 0 4224 0 1 15 0 0 2
221 211
181 211
1 4 4 0 0 8320 0 2 14 0 0 3
31 331
31 330
70 330
4 0 5 0 0 8320 0 5 0 0 26 4
386 451
385 451
385 193
218 193
17 4 5 0 0 0 0 13 5 0 0 3
418 459
418 451
386 451
3 18 6 0 0 8192 0 5 13 0 0 4
341 460
341 531
418 531
418 529
2 2 7 0 0 12416 0 4 5 0 0 6
422 348
421 348
421 343
311 343
311 451
341 451
2 3 6 0 0 8320 0 6 5 0 0 5
421 397
421 393
324 393
324 460
341 460
2 1 8 0 0 12416 0 3 5 0 0 5
421 306
421 300
303 300
303 442
341 442
1 0 9 0 0 4224 0 3 0 0 0 2
421 336
421 347
1 2 6 0 0 0 0 4 6 0 0 3
422 378
421 378
421 397
1 8 10 0 0 8320 0 6 12 0 0 3
421 433
421 434
448 434
1 19 2 0 0 12416 0 11 11 0 0 5
160 285
159 285
159 255
230 255
230 285
1 0 11 0 0 8192 0 19 0 0 17 4
151 604
151 539
253 539
253 540
2 0 12 0 0 8192 0 19 0 0 18 3
160 604
160 546
242 546
3 0 13 0 0 8192 0 19 0 0 19 3
169 604
169 554
233 554
4 0 14 0 0 8192 0 19 0 0 20 3
178 604
178 561
222 561
15 10 11 0 0 8320 0 11 13 0 0 5
224 339
253 339
253 540
436 540
436 529
16 12 12 0 0 12416 0 11 13 0 0 5
224 348
242 348
242 546
454 546
454 529
17 14 13 0 0 12416 0 11 13 0 0 5
224 357
233 357
233 554
472 554
472 529
18 16 14 0 0 12416 0 11 13 0 0 5
224 366
222 366
222 561
490 561
490 529
13 20 15 0 0 12416 0 15 11 0 0 6
117 157
112 157
112 249
242 249
242 294
230 294
1 11 16 0 0 12416 0 14 15 0 0 5
70 303
70 269
101 269
101 193
117 193
1 6 17 0 0 8320 0 8 15 0 0 5
64 243
64 242
195 242
195 166
181 166
3 1 17 0 0 0 0 14 8 0 0 2
64 321
64 243
3 2 17 0 0 0 0 14 14 0 0 3
64 321
64 312
70 312
7 3 5 0 0 0 0 15 15 0 0 4
181 157
218 157
218 193
181 193
3 2 18 0 0 4224 0 16 15 0 0 4
93 89
206 89
206 202
181 202
1 10 2 0 0 0 0 7 15 0 0 2
187 130
187 130
1 1 2 0 0 0 0 11 10 0 0 2
160 285
145 285
6 5 2 0 0 0 0 11 11 0 0 2
160 330
160 321
5 4 2 0 0 0 0 11 11 0 0 2
160 321
160 312
4 3 2 0 0 0 0 11 11 0 0 2
160 312
160 303
3 2 2 0 0 0 0 11 11 0 0 2
160 303
160 294
1 2 2 0 0 0 0 11 11 0 0 2
160 285
160 294
1 5 2 0 0 0 0 9 14 0 0 3
64 374
64 339
70 339
1 6 2 0 0 0 0 9 14 0 0 3
64 374
64 348
70 348
1 7 2 0 0 0 0 9 14 0 0 3
64 374
64 357
70 357
1 8 2 0 0 0 0 9 14 0 0 3
64 374
64 366
70 366
4 2 19 0 0 8320 0 12 13 0 0 4
472 434
472 442
436 442
436 465
3 4 20 0 0 8320 0 12 13 0 0 4
478 434
478 450
454 450
454 465
2 6 21 0 0 4224 0 12 13 0 0 4
484 434
484 457
472 457
472 465
8 1 22 0 0 4224 0 13 12 0 0 2
490 465
490 434
10 14 23 0 0 4224 0 11 14 0 0 2
160 366
134 366
9 13 24 0 0 4224 0 11 14 0 0 2
160 357
134 357
8 12 25 0 0 4224 0 11 14 0 0 2
160 348
134 348
7 11 26 0 0 4224 0 11 14 0 0 2
160 339
134 339
1 2 27 0 0 0 0 18 20 0 0 2
68 569
68 569
1 9 28 0 0 4224 0 20 17 0 0 2
68 605
68 604
1 13 29 0 0 8320 0 17 19 0 0 4
47 676
47 685
205 685
205 674
12 2 30 0 0 8320 0 19 17 0 0 4
196 674
196 684
53 684
53 676
11 3 31 0 0 8320 0 19 17 0 0 4
187 674
187 684
59 684
59 676
10 4 32 0 0 8320 0 19 17 0 0 4
178 674
178 684
65 684
65 676
8 6 33 0 0 8320 0 19 17 0 0 4
160 674
160 684
77 684
77 676
9 5 34 0 0 8320 0 19 17 0 0 4
169 674
169 684
71 684
71 676
7 7 35 0 0 8320 0 19 17 0 0 4
151 674
151 684
83 684
83 676
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 159
481 187 804 324
494 197 809 302
159 roll number dsiplay using counter and logic 
gates:

E (N) will be displayed by symbol display of 
14
and last letter will be blank (?)and then 
reset
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
