CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 1 80 9
0 70 1280 679
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1280 679
143654930 0
0
6 Title:
5 Name:
0
0
0
40
2 +V
167 298 575 0 1 3
0 8
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V4
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 617 584 0 1 3
0 7
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V2
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 74LS273
150 197 590 0 18 37
0 8 9 83 84 85 86 3 4 5
6 87 88 89 90 58 59 60 61
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U9
66 0 80 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3618 0 0
0
0
6 74LS47
187 708 1007 0 14 29
0 13 14 15 16 91 92 17 18 19
20 21 22 23 93
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
3 U17
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
6 74LS47
187 708 888 0 14 29
0 27 26 25 24 94 95 28 29 30
31 32 33 34 96
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
3 U16
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
6 74LS47
187 701 773 0 14 29
0 11 12 36 35 97 98 37 38 39
40 41 42 43 99
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
3 U15
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
6 74LS47
187 678 556 0 14 29
0 3 4 5 6 7 10 51 52 53
54 55 56 57 10
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
3 U14
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
7 74LS273
150 196 925 0 18 37
0 8 9 100 101 102 103 27 26 25
24 104 105 106 107 13 14 15 16
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
3 U13
61 -1 82 7
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
7 74LS273
150 197 800 0 18 37
0 8 9 108 109 110 111 11 12 36
35 112 113 114 115 27 26 25 24
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U1
62 -6 76 2
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
2 +V
167 847 423 0 1 3
0 62
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
9 CA 7-Seg~
184 848 575 0 18 19
10 23 22 21 20 19 18 17 116 67
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-44 -43 -9 -35
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9325 0 0
0
0
9 CA 7-Seg~
184 914 572 0 18 19
10 34 33 32 31 30 29 28 117 66
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
-47 -50 -12 -42
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8903 0 0
0
0
9 CA 7-Seg~
184 981 570 0 18 19
10 43 42 41 40 39 38 37 118 65
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
-46 -46 -11 -38
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3834 0 0
0
0
9 CA 7-Seg~
184 1041 569 0 18 19
10 50 49 48 47 46 45 44 119 64
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
-47 -43 -12 -35
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
9 CA 7-Seg~
184 1106 568 0 18 19
10 57 56 55 54 53 52 51 120 63
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
-47 -43 -12 -35
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7668 0 0
0
0
7 74LS273
150 196 707 0 18 37
0 8 9 121 122 123 124 58 59 60
61 125 126 127 128 11 12 36 35
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
3 U12
63 0 84 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
6 74LS47
187 760 671 0 14 29
0 58 59 60 61 129 130 44 45 46
47 48 49 50 131
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
3 U11
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
9 2-In AND~
219 113 466 0 3 22
0 68 69 70
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7C
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 5 0
1 U
6671 0 0
0
0
8 2-In OR~
219 71 504 0 3 22
0 70 71 4
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U8A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2010083361
65 0 0 0 4 1 6 0
1 U
3789 0 0
0
0
9 2-In AND~
219 43 344 0 3 22
0 68 73 72
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7B
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
4871 0 0
0
0
9 2-In AND~
219 67 299 0 3 22
0 74 73 71
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7A
4 13 25 21
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
3750 0 0
0
0
8 3-In OR~
219 23 457 0 4 22
0 71 72 69 3
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U6C
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 4 0
1 U
8778 0 0
0
0
9 2-In AND~
219 107 299 0 3 22
0 68 69 75
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4D
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
538 0 0
0
0
9 2-In AND~
219 146 299 0 3 22
0 74 68 76
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4C
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6843 0 0
0
0
8 3-In OR~
219 178 459 0 4 22
0 71 76 75 5
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U6B
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 4 0
1 U
3136 0 0
0
0
8 3-In OR~
219 224 424 0 4 22
0 77 78 79 6
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U6A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
5950 0 0
0
0
9 3-In AND~
219 177 346 0 4 22
0 80 74 68 79
0
0 0 624 270
6 74LS11
-21 -28 21 -20
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
5670 0 0
0
0
9 2-In AND~
219 230 349 0 3 22
0 81 82 78
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
6828 0 0
0
0
9 2-In AND~
219 285 347 0 3 22
0 73 81 77
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2093969452
65 0 0 0 4 1 2 0
1 U
6735 0 0
0
0
9 Inverter~
13 303 240 0 2 22
0 80 73
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
8365 0 0
0
0
9 Inverter~
13 256 239 0 2 22
0 74 81
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
4132 0 0
0
0
9 Inverter~
13 202 240 0 2 22
0 68 82
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
4551 0 0
0
0
7 Pulser~
4 69 98 0 10 12
0 132 133 10 9 0 0 5 5 6
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3635 0 0
0
0
6 74LS90
107 182 145 0 10 21
0 2 134 135 2 10 68 69 80 74
68
0
0 0 13040 270
6 74LS90
-21 -51 21 -43
2 U2
40 -4 54 4
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3973 0 0
0
0
7 Ground~
168 175 91 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3851 0 0
0
0
9 Resistor~
219 847 511 0 4 5
0 67 62 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 913 508 0 4 5
0 66 62 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 980 506 0 4 5
0 65 62 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 1040 505 0 4 5
0 64 62 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 1105 504 0 4 5
0 63 62 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
142
0 1 3 0 0 4240 0 0 7 8 0 2
26 520
646 520
2 0 4 0 0 4224 0 7 0 0 7 4
646 529
100 529
100 537
74 537
3 0 5 0 0 4224 0 7 0 0 6 2
646 538
181 538
4 0 6 0 0 4224 0 7 0 0 5 2
646 547
227 547
4 10 6 0 0 0 0 26 3 0 0 4
227 454
227 549
151 549
151 563
4 9 5 0 0 0 0 25 3 0 0 4
181 489
181 549
160 549
160 563
3 8 4 0 0 0 0 19 3 0 0 4
74 534
74 549
169 549
169 563
4 7 3 0 0 0 0 22 3 0 0 4
26 487
26 549
178 549
178 563
1 5 7 0 0 8320 0 2 7 0 0 3
617 593
617 592
646 592
1 0 8 0 0 4096 0 3 0 0 76 2
232 557
232 555
4 2 9 0 0 8320 0 33 3 0 0 5
99 98
341 98
341 543
223 543
223 563
3 6 10 0 0 8320 0 33 7 0 0 4
93 89
474 89
474 601
646 601
6 14 10 0 0 0 0 7 7 0 0 6
646 601
642 601
642 616
724 616
724 601
710 601
1 15 11 0 0 4224 0 6 16 0 0 5
669 737
250 737
250 711
177 711
177 744
2 0 12 0 0 8320 0 6 0 0 92 5
669 746
669 749
250 749
250 750
168 750
3 5 10 0 0 0 0 33 34 0 0 4
93 89
93 69
157 69
157 108
15 1 13 0 0 8320 0 8 4 0 0 3
177 962
177 971
676 971
16 2 14 0 0 8320 0 8 4 0 0 3
168 962
168 980
676 980
17 3 15 0 0 8320 0 8 4 0 0 3
159 962
159 989
676 989
18 4 16 0 0 8320 0 8 4 0 0 3
150 962
150 998
676 998
7 7 17 0 0 8320 0 4 11 0 0 3
746 971
863 971
863 611
8 6 18 0 0 8320 0 4 11 0 0 3
746 980
857 980
857 611
9 5 19 0 0 8320 0 4 11 0 0 3
746 989
851 989
851 611
10 4 20 0 0 8320 0 4 11 0 0 3
746 998
845 998
845 611
11 3 21 0 0 8320 0 4 11 0 0 3
746 1007
839 1007
839 611
12 2 22 0 0 8320 0 4 11 0 0 3
746 1016
833 1016
833 611
13 1 23 0 0 8320 0 4 11 0 0 3
746 1025
827 1025
827 611
4 0 24 0 0 4224 0 5 0 0 90 5
676 879
251 879
251 882
151 882
151 839
3 17 25 0 0 4224 0 5 9 0 0 5
676 870
251 870
251 873
160 873
160 837
2 0 26 0 0 4224 0 5 0 0 88 5
676 861
251 861
251 862
169 862
169 837
1 15 27 0 0 4224 0 5 9 0 0 5
676 852
251 852
251 855
178 855
178 837
7 0 28 0 0 4096 0 12 0 0 39 2
929 608
928 608
6 0 29 0 0 4096 0 12 0 0 40 2
923 608
922 608
5 0 30 0 0 4096 0 12 0 0 41 2
917 608
916 608
4 0 31 0 0 4096 0 12 0 0 42 2
911 608
910 608
3 0 32 0 0 4096 0 12 0 0 43 2
905 608
904 608
2 0 33 0 0 4096 0 12 0 0 44 2
899 608
898 608
1 0 34 0 0 4096 0 12 0 0 45 2
893 608
892 608
7 7 28 0 0 8320 0 5 0 0 0 3
746 852
928 852
928 604
8 6 29 0 0 8320 0 5 0 0 0 3
746 861
922 861
922 604
9 5 30 0 0 8320 0 5 0 0 0 3
746 870
916 870
916 604
10 4 31 0 0 8320 0 5 0 0 0 3
746 879
910 879
910 604
11 3 32 0 0 8320 0 5 0 0 0 3
746 888
904 888
904 604
12 2 33 0 0 8320 0 5 0 0 0 3
746 897
898 897
898 604
13 1 34 0 0 8320 0 5 0 0 0 3
746 906
892 906
892 604
4 18 35 0 0 8320 0 6 16 0 0 4
669 764
669 763
150 763
150 744
3 17 36 0 0 4224 0 6 16 0 0 3
669 755
159 755
159 744
7 0 37 0 0 0 0 13 0 0 55 2
996 606
996 606
6 0 38 0 0 0 0 13 0 0 56 2
990 606
990 606
5 0 39 0 0 0 0 13 0 0 57 2
984 606
984 606
4 0 40 0 0 0 0 13 0 0 58 2
978 606
978 606
3 0 41 0 0 0 0 13 0 0 59 2
972 606
972 606
2 0 42 0 0 0 0 13 0 0 60 2
966 606
966 606
1 0 43 0 0 0 0 13 0 0 61 2
960 606
960 606
7 7 37 0 0 4224 0 6 0 0 0 3
739 737
996 737
996 602
8 6 38 0 0 4224 0 6 0 0 0 3
739 746
990 746
990 602
9 5 39 0 0 4224 0 6 0 0 0 3
739 755
984 755
984 602
10 4 40 0 0 4224 0 6 0 0 0 3
739 764
978 764
978 602
11 3 41 0 0 4224 0 6 0 0 0 3
739 773
972 773
972 602
12 2 42 0 0 4224 0 6 0 0 0 3
739 782
966 782
966 602
13 1 43 0 0 4224 0 6 0 0 0 3
739 791
960 791
960 602
7 7 44 0 0 4224 0 17 14 0 0 3
798 635
1056 635
1056 605
8 6 45 0 0 4224 0 17 14 0 0 3
798 644
1050 644
1050 605
9 5 46 0 0 4224 0 17 14 0 0 3
798 653
1044 653
1044 605
10 4 47 0 0 4224 0 17 14 0 0 3
798 662
1038 662
1038 605
11 3 48 0 0 4224 0 17 14 0 0 3
798 671
1032 671
1032 605
12 2 49 0 0 4224 0 17 14 0 0 3
798 680
1026 680
1026 605
13 1 50 0 0 4224 0 17 14 0 0 3
798 689
1020 689
1020 605
7 7 51 0 0 12416 0 7 15 0 0 5
716 520
818 520
818 616
1121 616
1121 604
8 6 52 0 0 12416 0 7 15 0 0 5
716 529
818 529
818 616
1115 616
1115 604
9 5 53 0 0 12416 0 7 15 0 0 5
716 538
818 538
818 616
1109 616
1109 604
10 4 54 0 0 12416 0 7 15 0 0 5
716 547
818 547
818 616
1103 616
1103 604
11 3 55 0 0 12416 0 7 15 0 0 5
716 556
818 556
818 616
1097 616
1097 604
12 2 56 0 0 12416 0 7 15 0 0 5
716 565
818 565
818 616
1091 616
1091 604
13 1 57 0 0 12416 0 7 15 0 0 5
716 574
818 574
818 616
1085 616
1085 604
1 0 8 0 0 20480 0 1 0 0 10 7
298 584
285 584
285 561
286 561
286 555
232 555
232 557
0 1 58 0 0 4224 0 0 17 95 0 2
178 635
728 635
0 2 59 0 0 4224 0 0 17 96 0 2
169 644
728 644
0 3 60 0 0 4224 0 0 17 97 0 3
160 654
728 654
728 653
0 4 61 0 0 4224 0 0 17 98 0 3
151 663
728 663
728 662
0 2 9 0 0 0 0 0 8 82 0 4
341 770
341 835
222 835
222 898
0 2 9 0 0 0 0 0 9 83 0 5
342 669
341 669
341 770
223 770
223 773
0 2 9 0 0 0 0 0 16 11 0 7
341 543
343 543
343 595
342 595
342 670
222 670
222 680
0 1 8 0 0 4096 0 0 8 85 0 4
274 766
274 840
231 840
231 892
0 1 8 0 0 4096 0 0 9 86 0 4
274 674
274 766
232 766
232 767
0 1 8 0 0 16512 0 0 16 76 0 6
285 561
284 561
284 556
274 556
274 674
231 674
7 15 27 0 0 0 0 8 9 0 0 4
177 898
177 840
178 840
178 837
8 16 26 0 0 0 0 8 9 0 0 3
168 898
168 837
169 837
9 17 25 0 0 0 0 8 9 0 0 4
159 898
159 840
160 840
160 837
10 18 24 0 0 0 0 8 9 0 0 4
150 898
150 839
151 839
151 837
7 15 11 0 0 0 0 9 16 0 0 4
178 773
178 762
177 762
177 744
8 16 12 0 0 0 0 9 16 0 0 4
169 773
169 754
168 754
168 744
9 17 36 0 0 0 0 9 16 0 0 4
160 773
160 762
159 762
159 744
10 18 35 0 0 0 0 9 16 0 0 4
151 773
151 762
150 762
150 744
7 15 58 0 0 0 0 16 3 0 0 4
177 680
177 635
178 635
178 627
8 16 59 0 0 0 0 16 3 0 0 4
168 680
168 644
169 644
169 627
9 17 60 0 0 0 0 16 3 0 0 4
159 680
159 654
160 654
160 627
10 18 61 0 0 0 0 16 3 0 0 4
150 680
150 663
151 663
151 627
1 2 62 0 0 8320 0 10 40 0 0 4
847 432
847 478
1105 478
1105 486
1 2 62 0 0 0 0 10 39 0 0 4
847 432
847 462
1040 462
1040 487
1 2 62 0 0 0 0 10 38 0 0 5
847 432
846 432
846 454
980 454
980 488
1 2 62 0 0 0 0 10 37 0 0 4
847 432
847 442
913 442
913 490
1 9 63 0 0 8320 0 40 15 0 0 3
1105 522
1106 522
1106 532
1 9 64 0 0 8320 0 39 14 0 0 3
1040 523
1041 523
1041 533
1 9 65 0 0 8320 0 38 13 0 0 3
980 524
981 524
981 534
1 9 66 0 0 8320 0 37 12 0 0 3
913 526
914 526
914 536
1 2 62 0 0 0 0 10 36 0 0 2
847 432
847 493
1 9 67 0 0 8320 0 36 11 0 0 3
847 529
848 529
848 539
1 1 68 0 0 4096 0 18 20 0 0 4
120 444
120 347
50 347
50 322
2 0 69 0 0 12288 0 18 0 0 120 4
102 444
97 444
97 396
17 396
3 1 70 0 0 8320 0 18 19 0 0 4
111 489
111 487
83 487
83 488
2 0 71 0 0 4096 0 19 0 0 116 2
65 488
65 420
1 0 68 0 0 0 0 20 0 0 122 4
50 322
45 322
45 258
114 258
3 2 72 0 0 8320 0 20 22 0 0 3
41 367
26 367
26 442
2 0 73 0 0 4096 0 20 0 0 118 3
32 322
32 266
56 266
1 0 71 0 0 0 0 22 0 0 119 3
35 441
35 420
65 420
1 0 74 0 0 8192 0 21 0 0 126 3
74 277
74 248
158 248
2 0 73 0 0 8320 0 21 0 0 135 3
56 277
56 266
306 266
3 1 71 0 0 8320 0 21 25 0 0 4
65 322
65 420
190 420
190 443
3 0 69 0 0 4224 0 22 0 0 121 3
17 441
17 232
96 232
2 7 69 0 0 0 0 23 34 0 0 4
96 277
96 184
202 184
202 178
1 0 68 0 0 0 0 23 0 0 125 3
114 277
114 257
135 257
3 3 75 0 0 4224 0 23 25 0 0 4
105 322
105 437
172 437
172 443
3 2 76 0 0 4224 0 24 25 0 0 4
144 322
144 428
181 428
181 444
2 0 68 0 0 0 0 24 0 0 139 3
135 277
135 200
148 200
1 0 74 0 0 0 0 24 0 0 138 4
153 277
158 277
158 199
166 199
1 3 77 0 0 8320 0 26 29 0 0 4
236 408
236 378
283 378
283 370
2 3 78 0 0 4224 0 26 28 0 0 4
227 409
227 380
228 380
228 372
3 4 79 0 0 8320 0 26 27 0 0 4
218 408
218 376
175 376
175 369
1 0 80 0 0 4224 0 27 0 0 137 2
184 324
184 189
2 0 74 0 0 4224 0 27 0 0 138 2
175 324
175 201
3 0 68 0 0 4224 0 27 0 0 139 2
166 324
166 214
2 1 81 0 0 8320 0 31 28 0 0 5
259 257
255 257
255 319
237 319
237 327
2 2 82 0 0 4224 0 32 28 0 0 4
205 258
205 319
219 319
219 327
2 1 73 0 0 0 0 30 29 0 0 4
306 258
306 317
292 317
292 325
2 2 81 0 0 0 0 31 29 0 0 5
259 257
262 257
262 317
274 317
274 325
8 1 80 0 0 0 0 34 30 0 0 4
184 178
184 189
306 189
306 222
9 1 74 0 0 0 0 34 31 0 0 4
166 178
166 201
259 201
259 221
10 1 68 0 0 0 0 34 32 0 0 4
148 178
148 214
205 214
205 222
1 0 2 0 0 0 0 35 0 0 141 2
175 99
175 99
4 1 2 0 0 8320 0 34 34 0 0 4
175 114
175 99
202 99
202 114
6 10 68 0 0 0 0 34 34 0 0 6
148 108
148 103
134 103
134 177
148 177
148 178
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
