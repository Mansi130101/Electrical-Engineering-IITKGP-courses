CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 E:\CircuitMaker\BOM.DAT
0 7
0 71 1536 824
143654930 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 518 349 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
7 Pulser~
4 443 94 0 10 12
0 50 51 3 52 0 0 5 5 5
8
0
0 0 4656 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4441 0 0
0
0
7 Pulser~
4 111 91 0 10 12
0 53 54 2 55 0 0 5 5 5
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3618 0 0
0
0
2 +V
167 265 63 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
2 +V
167 539 61 0 1 3
0 5
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
2 +V
167 1128 285 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
2 +V
167 982 279 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
7 74LS273
150 593 146 0 18 37
0 5 3 34 35 36 37 38 39 40
41 26 27 28 29 30 31 32 33
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
7 74LS273
150 321 146 0 18 37
0 4 2 45 44 43 42 46 47 48
49 34 35 36 37 38 39 40 41
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
6 74LS83
105 400 351 0 14 29
0 33 32 31 30 41 40 39 38 25
49 48 47 46 56
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
6 74LS83
105 620 354 0 14 29
0 29 28 27 26 37 36 35 34 24
42 43 44 45 25
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U3
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
6 74LS47
187 838 639 0 14 29
0 42 43 44 45 57 58 10 11 12
13 14 15 16 59
0
0 0 13040 0
7 74LS247
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
6 74LS47
187 839 512 0 14 29
0 49 48 47 46 60 61 17 18 19
20 21 22 23 62
0
0 0 13040 0
7 74LS247
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
9 CA 7-Seg~
184 1128 395 0 18 19
10 16 15 14 13 12 11 10 63 9
0 0 0 2 2 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3363 0 0
0
0
9 CA 7-Seg~
184 982 394 0 18 19
10 23 22 21 20 19 18 17 64 7
2 2 2 0 0 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7668 0 0
0
0
9 Resistor~
219 1128 325 0 4 5
0 9 8 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 982 321 0 4 5
0 7 6 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3874 0 0
0
0
64
3 2 2 0 0 4224 0 3 9 0 0 4
135 82
251 82
251 119
289 119
3 2 3 0 0 4224 0 2 8 0 0 4
467 85
526 85
526 119
561 119
1 1 4 0 0 8320 0 9 4 0 0 3
283 110
265 110
265 72
1 1 5 0 0 4224 0 5 8 0 0 3
539 70
539 110
555 110
2 1 6 0 0 4224 0 17 7 0 0 2
982 303
982 288
9 1 7 0 0 4224 0 15 17 0 0 2
982 358
982 339
2 1 8 0 0 4224 0 16 6 0 0 2
1128 307
1128 294
9 1 9 0 0 4224 0 14 16 0 0 2
1128 359
1128 343
7 7 10 0 0 4224 0 12 14 0 0 3
876 603
1143 603
1143 431
8 6 11 0 0 4224 0 12 14 0 0 3
876 612
1137 612
1137 431
9 5 12 0 0 4224 0 12 14 0 0 3
876 621
1131 621
1131 431
10 4 13 0 0 4224 0 12 14 0 0 3
876 630
1125 630
1125 431
11 3 14 0 0 4224 0 12 14 0 0 3
876 639
1119 639
1119 431
12 2 15 0 0 4224 0 12 14 0 0 3
876 648
1113 648
1113 431
13 1 16 0 0 4224 0 12 14 0 0 3
876 657
1107 657
1107 431
7 7 17 0 0 4224 0 13 15 0 0 3
877 476
997 476
997 430
8 6 18 0 0 4224 0 13 15 0 0 3
877 485
991 485
991 430
9 5 19 0 0 4224 0 13 15 0 0 3
877 494
985 494
985 430
10 4 20 0 0 4224 0 13 15 0 0 3
877 503
979 503
979 430
11 3 21 0 0 4224 0 13 15 0 0 3
877 512
973 512
973 430
12 2 22 0 0 8320 0 13 15 0 0 3
877 521
967 521
967 430
13 1 23 0 0 8320 0 13 15 0 0 3
877 530
961 530
961 430
1 9 24 0 0 8320 0 1 11 0 0 5
530 349
552 349
552 311
577 311
577 324
14 9 25 0 0 8320 0 11 10 0 0 6
577 388
577 397
331 397
331 299
357 299
357 321
4 11 26 0 0 12416 0 11 8 0 0 5
631 324
631 302
731 302
731 128
625 128
12 3 27 0 0 8320 0 8 11 0 0 5
625 137
718 137
718 293
640 293
640 324
2 13 28 0 0 12416 0 11 8 0 0 5
649 324
649 286
706 286
706 146
625 146
14 1 29 0 0 8320 0 8 11 0 0 5
625 155
694 155
694 277
658 277
658 324
15 4 30 0 0 12416 0 8 10 0 0 5
625 164
685 164
685 246
411 246
411 321
3 16 31 0 0 8320 0 10 8 0 0 5
420 321
420 234
674 234
674 173
625 173
17 2 32 0 0 12416 0 8 10 0 0 5
625 182
663 182
663 224
429 224
429 321
1 18 33 0 0 8320 0 10 8 0 0 5
438 321
438 211
653 211
653 191
625 191
8 0 34 0 0 12288 0 11 0 0 57 4
595 324
595 303
499 303
499 128
7 0 35 0 0 12288 0 11 0 0 58 4
604 324
604 293
510 293
510 137
6 0 36 0 0 12288 0 11 0 0 59 4
613 324
613 284
520 284
520 146
5 0 37 0 0 12288 0 11 0 0 60 4
622 324
622 276
529 276
529 155
8 0 38 0 0 4096 0 10 0 0 61 2
375 321
375 164
7 0 39 0 0 4096 0 10 0 0 62 2
384 321
384 173
6 0 40 0 0 4096 0 10 0 0 63 2
393 321
393 182
5 0 41 0 0 4096 0 10 0 0 64 2
402 321
402 191
6 0 42 0 0 12416 0 9 0 0 49 4
289 155
192 155
192 573
631 573
5 0 43 0 0 12416 0 9 0 0 50 4
289 146
180 146
180 563
622 563
4 0 44 0 0 12416 0 9 0 0 51 4
289 137
169 137
169 553
613 553
3 0 45 0 0 12416 0 9 0 0 52 4
289 128
160 128
160 543
604 543
7 0 46 0 0 8192 0 9 0 0 56 4
289 164
229 164
229 440
384 440
8 0 47 0 0 8192 0 9 0 0 55 4
289 173
240 173
240 428
393 428
9 0 48 0 0 8192 0 9 0 0 54 4
289 182
249 182
249 419
402 419
10 0 49 0 0 8192 0 9 0 0 53 4
289 191
258 191
258 410
411 410
10 1 42 0 0 0 0 11 12 0 0 3
631 388
631 603
806 603
11 2 43 0 0 0 0 11 12 0 0 3
622 388
622 612
806 612
12 3 44 0 0 0 0 11 12 0 0 3
613 388
613 621
806 621
13 4 45 0 0 0 0 11 12 0 0 3
604 388
604 630
806 630
10 1 49 0 0 8320 0 10 13 0 0 3
411 385
411 476
807 476
2 11 48 0 0 4224 0 13 10 0 0 3
807 485
402 485
402 385
12 3 47 0 0 8320 0 10 13 0 0 3
393 385
393 494
807 494
13 4 46 0 0 8320 0 10 13 0 0 3
384 385
384 503
807 503
11 3 34 0 0 4224 0 9 8 0 0 2
353 128
561 128
12 4 35 0 0 4224 0 9 8 0 0 2
353 137
561 137
13 5 36 0 0 4224 0 9 8 0 0 2
353 146
561 146
14 6 37 0 0 4224 0 9 8 0 0 2
353 155
561 155
15 7 38 0 0 4224 0 9 8 0 0 2
353 164
561 164
16 8 39 0 0 4224 0 9 8 0 0 2
353 173
561 173
17 9 40 0 0 4224 0 9 8 0 0 2
353 182
561 182
18 10 41 0 0 4224 0 9 8 0 0 2
353 191
561 191
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
