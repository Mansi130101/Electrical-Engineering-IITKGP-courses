CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 25 100 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
143654930 0
0
6 Title:
5 Name:
0
0
0
26
9 CA 7-Seg~
184 806 158 0 18 19
10 14 13 12 11 10 9 8 58 16
0 2 0 0 2 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8953 0 0
0
0
2 +V
167 806 61 0 1 3
0 15
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
6 74LS47
187 794 253 0 14 29
0 3 7 4 5 59 60 8 9 10
11 12 13 14 61
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U6
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3618 0 0
0
0
6 74LS93
109 828 335 0 8 17
0 3 4 6 5 3 7 4 5
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U5
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
7 Pulser~
4 735 391 0 10 12
0 62 63 6 64 0 0 5 5 1
7
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5394 0 0
0
0
9 2-In AND~
219 375 489 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
4 15 25 23
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 800149019
65 0 0 0 4 3 1 0
1 U
7734 0 0
0
0
8 2-In OR~
219 407 435 0 3 22
0 22 19 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 565267989
65 0 0 0 4 1 2 0
1 U
9914 0 0
0
0
9 2-In AND~
219 273 253 0 3 22
0 17 23 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 800149019
65 0 0 0 4 2 1 0
1 U
3747 0 0
0
0
9 2-In AND~
219 280 415 0 3 22
0 17 23 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 615599632
65 0 0 0 4 1 1 0
1 U
3549 0 0
0
0
7 Ground~
168 189 257 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
6 74LS93
109 147 311 0 8 17
0 24 65 19 25 17 17 17 25
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U8
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
6 74LS47
187 113 229 0 14 29
0 2 2 17 25 66 67 26 27 28
29 30 31 32 68
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
2 +V
167 125 37 0 1 3
0 33
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
9 CA 7-Seg~
184 125 129 0 18 19
10 32 31 30 29 28 27 26 69 34
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
9 CA 7-Seg~
184 416 145 0 18 19
10 43 42 41 40 39 38 37 70 45
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7668 0 0
0
0
2 +V
167 416 48 0 1 3
0 44
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
6 74LS47
187 404 240 0 14 29
0 21 23 20 36 71 72 37 38 39
40 41 42 43 73
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
6 74LS93
109 438 322 0 8 17
0 18 74 35 36 21 23 20 36
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U3
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
9 CA 7-Seg~
184 578 159 0 18 19
10 55 54 53 52 51 50 49 75 57
0 0 0 0 2 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3789 0 0
0
0
2 +V
167 578 62 0 1 3
0 56
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4871 0 0
0
0
6 74LS47
187 566 254 0 14 29
0 48 35 46 47 76 77 49 50 51
52 53 54 55 78
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
6 74LS93
109 600 336 0 8 17
0 35 46 3 47 48 35 46 47
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U1
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
9 Resistor~
219 806 96 0 4 5
0 16 15 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 125 72 0 4 5
0 34 33 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 416 83 0 4 5
0 45 44 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 578 97 0 4 5
0 57 56 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
76
3 0 3 0 0 8320 0 22 0 0 3 4
589 372
589 420
861 420
861 373
2 0 4 0 0 12416 0 4 0 0 7 5
826 365
826 381
887 381
887 294
817 294
1 5 3 0 0 0 0 4 4 0 0 5
835 365
835 373
875 373
875 301
835 301
4 0 5 0 0 12416 0 4 0 0 6 5
808 371
808 375
793 375
793 301
808 301
3 3 6 0 0 4224 0 5 4 0 0 4
759 382
816 382
816 371
817 371
8 4 5 0 0 0 0 4 3 0 0 2
808 301
808 290
7 3 4 0 0 0 0 4 3 0 0 2
817 301
817 290
6 2 7 0 0 4224 0 4 3 0 0 2
826 301
826 290
5 1 3 0 0 0 0 4 3 0 0 2
835 301
835 290
7 7 8 0 0 4224 0 3 1 0 0 4
835 220
835 200
821 200
821 194
8 6 9 0 0 4224 0 3 1 0 0 4
826 220
826 203
815 203
815 194
9 5 10 0 0 12416 0 3 1 0 0 4
817 220
817 208
809 208
809 194
10 4 11 0 0 12416 0 3 1 0 0 4
808 220
808 213
803 213
803 194
11 3 12 0 0 4224 0 3 1 0 0 4
799 220
799 202
797 202
797 194
12 2 13 0 0 4224 0 3 1 0 0 4
790 220
790 201
791 201
791 194
13 1 14 0 0 4224 0 3 1 0 0 4
781 220
781 202
785 202
785 194
1 2 15 0 0 4224 0 2 23 0 0 2
806 70
806 78
1 9 16 0 0 4224 0 23 1 0 0 2
806 114
806 122
1 2 2 0 0 4096 0 12 12 0 0 2
154 266
145 266
1 1 2 0 0 12416 0 10 12 0 0 5
189 251
189 247
173 247
173 266
154 266
6 0 17 0 0 0 0 11 0 0 33 2
145 277
145 277
5 0 17 0 0 0 0 11 0 0 33 2
154 277
154 277
3 1 18 0 0 8320 0 7 18 0 0 3
440 435
445 435
445 352
3 0 19 0 0 8320 0 11 0 0 27 3
136 347
136 465
394 465
2 7 20 0 0 16512 0 6 18 0 0 6
351 498
340 498
340 517
474 517
474 288
427 288
1 1 21 0 0 16512 0 6 17 0 0 6
351 480
319 480
319 527
496 527
496 277
445 277
3 2 19 0 0 0 0 6 7 0 0 3
396 489
394 489
394 444
3 1 22 0 0 8320 0 8 7 0 0 4
294 253
316 253
316 426
394 426
0 2 23 0 0 4096 0 0 8 32 0 4
338 282
245 282
245 262
249 262
0 1 17 0 0 4096 0 0 8 33 0 3
231 277
231 244
249 244
1 3 24 0 0 8320 0 11 9 0 0 4
154 341
154 355
301 355
301 415
2 2 23 0 0 12432 0 17 9 0 0 7
436 277
436 281
338 281
338 448
240 448
240 424
256 424
7 1 17 0 0 8320 0 11 9 0 0 4
136 277
231 277
231 406
256 406
4 0 25 0 0 12416 0 11 0 0 35 5
127 347
127 348
112 348
112 277
127 277
8 4 25 0 0 0 0 11 12 0 0 2
127 277
127 266
7 3 17 0 0 0 0 11 12 0 0 2
136 277
136 266
7 7 26 0 0 4224 0 12 14 0 0 4
154 196
154 176
140 176
140 165
8 6 27 0 0 4224 0 12 14 0 0 4
145 196
145 179
134 179
134 165
9 5 28 0 0 12416 0 12 14 0 0 4
136 196
136 184
128 184
128 165
10 4 29 0 0 12416 0 12 14 0 0 4
127 196
127 189
122 189
122 165
11 3 30 0 0 4224 0 12 14 0 0 4
118 196
118 178
116 178
116 165
12 2 31 0 0 4224 0 12 14 0 0 4
109 196
109 177
110 177
110 165
13 1 32 0 0 4224 0 12 14 0 0 4
100 196
100 178
104 178
104 165
1 2 33 0 0 4224 0 13 24 0 0 2
125 46
125 54
1 9 34 0 0 4224 0 24 14 0 0 4
125 90
125 94
125 94
125 93
0 3 35 0 0 12416 0 0 18 66 0 5
598 297
677 297
677 395
427 395
427 358
4 0 36 0 0 8320 0 18 0 0 48 4
418 358
403 358
403 288
418 288
8 4 36 0 0 0 0 18 17 0 0 2
418 288
418 277
7 3 20 0 0 0 0 18 17 0 0 2
427 288
427 277
6 2 23 0 0 0 0 18 17 0 0 2
436 288
436 277
5 1 21 0 0 0 0 18 17 0 0 2
445 288
445 277
7 7 37 0 0 4224 0 17 15 0 0 4
445 207
445 187
431 187
431 181
8 6 38 0 0 4224 0 17 15 0 0 4
436 207
436 190
425 190
425 181
9 5 39 0 0 12416 0 17 15 0 0 4
427 207
427 195
419 195
419 181
10 4 40 0 0 12416 0 17 15 0 0 4
418 207
418 200
413 200
413 181
11 3 41 0 0 4224 0 17 15 0 0 4
409 207
409 189
407 189
407 181
12 2 42 0 0 4224 0 17 15 0 0 4
400 207
400 188
401 188
401 181
13 1 43 0 0 4224 0 17 15 0 0 4
391 207
391 189
395 189
395 181
1 2 44 0 0 4224 0 16 25 0 0 2
416 57
416 65
1 9 45 0 0 4224 0 25 15 0 0 2
416 101
416 109
2 3 46 0 0 12416 0 22 21 0 0 5
598 366
598 379
653 379
653 291
589 291
1 6 35 0 0 0 0 22 22 0 0 5
607 366
607 373
645 373
645 302
598 302
4 0 47 0 0 12416 0 22 0 0 64 5
580 372
580 376
565 376
565 302
580 302
8 4 47 0 0 0 0 22 21 0 0 2
580 302
580 291
7 3 46 0 0 0 0 22 21 0 0 2
589 302
589 291
6 2 35 0 0 0 0 22 21 0 0 2
598 302
598 291
5 1 48 0 0 4224 0 22 21 0 0 2
607 302
607 291
7 7 49 0 0 4224 0 21 19 0 0 4
607 221
607 201
593 201
593 195
8 6 50 0 0 4224 0 21 19 0 0 4
598 221
598 204
587 204
587 195
9 5 51 0 0 12416 0 21 19 0 0 4
589 221
589 209
581 209
581 195
10 4 52 0 0 12416 0 21 19 0 0 4
580 221
580 214
575 214
575 195
11 3 53 0 0 4224 0 21 19 0 0 4
571 221
571 203
569 203
569 195
12 2 54 0 0 4224 0 21 19 0 0 4
562 221
562 202
563 202
563 195
13 1 55 0 0 4224 0 21 19 0 0 4
553 221
553 203
557 203
557 195
1 2 56 0 0 4224 0 20 26 0 0 2
578 71
578 79
1 9 57 0 0 4224 0 26 19 0 0 2
578 115
578 123
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
998 73 1110 117
1008 81 1112 113
25 MANSI UNIYAL 
19EE10039
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 704
932 124 1228 608
942 132 1230 516
704 For creating minutes display:

1. units place of minutes display 
would reset at 9 (ie. modulus 10).
2. tens place of minutes display 
would reset on 5 (ie. modulus 6) 
and take input when units place 
resets from 9 to 0. (as the maximum 
minutes is till 59)

For creating hours display:

1. units place of hours display 
would reset on 9 (ie. modulus 10)or 
when tens place displays 2 and 
units place displays 4.
2. units place of hours display 
takes input when tens place of 
minutes display resets from 5 to 0.
2. tens place of hours display 
takes input when units place of 
hours display resets from 9 to 0.
3. tens place of hours resets when 
hours display 24.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
