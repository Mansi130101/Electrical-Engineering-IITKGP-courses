CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 80 9
0 82 1920 1030
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 82 1920 1030
143654930 0
0
6 Title:
5 Name:
0
0
0
39
2 +V
167 947 254 0 1 3
0 4
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 890 39 0 1 3
0 5
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
9 CA 7-Seg~
184 249 97 0 18 19
10 17 16 15 14 13 12 11 84 10
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3618 0 0
0
0
9 CA 7-Seg~
184 394 97 0 18 19
10 24 23 22 21 20 19 18 85 9
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6153 0 0
0
0
9 CA 7-Seg~
184 531 96 0 18 19
10 31 30 29 28 27 26 25 86 8
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
9 CA 7-Seg~
184 664 99 0 18 19
10 38 37 36 35 34 33 32 87 7
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7734 0 0
0
0
9 CA 7-Seg~
184 794 99 0 18 19
10 45 44 43 42 41 40 39 88 6
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9914 0 0
0
0
6 74LS47
187 256 186 0 14 29
0 46 47 48 49 89 90 11 12 13
14 15 16 17 91
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
3 U17
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
6 74LS47
187 403 189 0 14 29
0 50 51 52 53 92 93 18 19 20
21 22 23 24 94
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
3 U16
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
6 74LS47
187 538 187 0 14 29
0 54 55 56 57 95 96 25 26 27
28 29 30 31 97
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
3 U15
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
6 74LS47
187 673 186 0 14 29
0 58 59 60 61 98 99 32 33 34
35 36 37 38 100
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
3 U14
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
6 74LS47
187 801 184 0 14 29
0 62 63 64 65 101 102 39 40 41
42 43 44 45 103
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
3 U13
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
7 Pulser~
4 1174 941 0 10 12
0 104 105 3 106 0 0 20 20 21
7
0
0 0 4656 512
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3834 0 0
0
0
6 74LS90
107 970 865 0 10 21
0 2 2 2 2 3 69 75 71 72
69
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U2
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
9 Inverter~
13 1025 738 0 2 22
0 69 73
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
7668 0 0
0
0
9 Inverter~
13 1071 739 0 2 22
0 72 78
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
4718 0 0
0
0
9 Inverter~
13 1117 741 0 2 22
0 71 68
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
3874 0 0
0
0
7 Ground~
168 984 914 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
5 4081~
219 949 642 0 3 22
0 72 68 79
0
0 0 624 90
4 4081
-7 -24 21 -16
3 U4A
16 -5 37 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3789 0 0
0
0
5 4081~
219 1017 641 0 3 22
0 69 75 83
0
0 0 624 90
4 4081
-7 -24 21 -16
3 U4B
16 -5 37 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
4871 0 0
0
0
5 4071~
219 981 482 0 3 22
0 79 83 82
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U5A
28 -3 49 5
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 3 0
1 U
3750 0 0
0
0
5 4071~
219 921 483 0 3 22
0 77 82 81
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U5B
28 -3 49 5
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 3 0
1 U
8778 0 0
0
0
8 3-In OR~
219 757 484 0 4 22
0 76 74 70 66
0
0 0 624 90
4 4075
-14 -24 14 -16
3 U6A
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
538 0 0
0
0
8 3-In OR~
219 1152 485 0 4 22
0 79 75 67 80
0
0 0 624 90
4 4075
-14 -24 14 -16
3 U6B
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 4 0
1 U
6843 0 0
0
0
5 4073~
219 898 560 0 4 22
0 73 78 71 77
0
0 0 624 90
4 4073
-7 -24 21 -16
3 U8A
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 6 0
1 U
3136 0 0
0
0
5 4073~
219 702 563 0 4 22
0 69 72 71 76
0
0 0 624 90
4 4073
-7 -24 21 -16
3 U8B
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 6 0
1 U
5950 0 0
0
0
5 4025~
219 754 562 0 4 22
0 69 72 75 74
0
0 0 624 90
4 4025
-14 -24 14 -16
3 U9A
31 0 52 8
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 7 0
1 U
5670 0 0
0
0
5 4025~
219 817 560 0 4 22
0 73 72 71 70
0
0 0 624 90
4 4025
-14 -24 14 -16
3 U9B
31 0 52 8
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 7 0
1 U
6828 0 0
0
0
5 4081~
219 1174 589 0 3 22
0 69 68 67
0
0 0 624 90
4 4081
-7 -24 21 -16
3 U4C
16 -5 37 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6735 0 0
0
0
7 74LS273
150 321 328 0 18 37
0 4 3 107 108 109 110 50 51 52
53 111 112 113 114 46 47 48 49
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
3 U12
-17 -61 4 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
8365 0 0
0
0
7 74LS273
150 450 330 0 18 37
0 4 3 115 116 117 118 54 55 56
57 119 120 121 122 50 51 52 53
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
3 U11
-17 -61 4 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
4132 0 0
0
0
7 74LS273
150 596 331 0 18 37
0 4 3 123 124 125 126 58 59 60
61 127 128 129 130 54 55 56 57
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
3 U10
-17 -61 4 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
4551 0 0
0
0
7 74LS273
150 721 332 0 18 37
0 4 3 131 132 133 134 62 63 64
65 135 136 137 138 58 59 60 61
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
2 U7
-13 -61 1 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3635 0 0
0
0
7 74LS273
150 840 333 0 18 37
0 4 3 139 140 141 142 80 82 81
66 143 144 145 146 62 63 64 65
0
0 0 13040 512
7 74LS273
-24 -60 25 -52
2 U1
-13 -61 1 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3973 0 0
0
0
9 Resistor~
219 249 34 0 4 5
0 10 5 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 393 33 0 4 5
0 9 5 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 531 36 0 4 5
0 8 5 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 664 35 0 4 5
0 7 5 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 793 34 0 4 5
0 6 5 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
132
2 0 3 0 0 8192 0 33 0 0 4 3
747 305
761 305
761 264
2 0 3 0 0 0 0 32 0 0 4 3
622 304
634 304
634 264
2 0 3 0 0 0 0 31 0 0 4 3
476 303
493 303
493 264
0 2 3 0 0 8320 0 0 30 5 0 5
913 306
913 264
361 264
361 301
347 301
2 0 3 0 0 0 0 34 0 0 128 5
866 306
1233 306
1233 801
1091 801
1091 932
1 0 4 0 0 4096 0 34 0 0 10 2
872 297
872 253
1 0 4 0 0 0 0 33 0 0 10 2
753 296
753 253
1 0 4 0 0 0 0 32 0 0 10 2
628 295
628 253
1 0 4 0 0 0 0 31 0 0 10 2
482 294
482 253
1 1 4 0 0 4224 0 1 30 0 0 3
935 253
353 253
353 292
2 0 5 0 0 4096 0 36 0 0 15 2
393 15
393 7
2 0 5 0 0 4096 0 37 0 0 15 2
531 18
531 7
2 0 5 0 0 0 0 38 0 0 15 2
664 17
664 7
2 0 5 0 0 0 0 39 0 0 15 2
793 16
793 7
2 1 5 0 0 8320 0 35 2 0 0 5
249 16
249 7
873 7
873 38
878 38
1 9 6 0 0 8320 0 39 7 0 0 3
793 52
794 52
794 63
1 9 7 0 0 4224 0 38 6 0 0 2
664 53
664 63
1 9 8 0 0 4224 0 37 5 0 0 2
531 54
531 60
1 9 9 0 0 8320 0 36 4 0 0 3
393 51
394 51
394 61
1 9 10 0 0 4224 0 35 3 0 0 2
249 52
249 61
7 7 11 0 0 8320 0 3 8 0 0 4
264 133
264 145
221 145
221 153
6 8 12 0 0 8320 0 3 8 0 0 4
258 133
258 145
230 145
230 153
5 9 13 0 0 8320 0 3 8 0 0 4
252 133
252 145
239 145
239 153
4 10 14 0 0 4224 0 3 8 0 0 4
246 133
246 145
248 145
248 153
3 11 15 0 0 8320 0 3 8 0 0 4
240 133
240 145
257 145
257 153
2 12 16 0 0 8320 0 3 8 0 0 4
234 133
234 145
266 145
266 153
1 13 17 0 0 8320 0 3 8 0 0 4
228 133
228 145
275 145
275 153
7 7 18 0 0 8320 0 4 9 0 0 4
409 133
409 148
368 148
368 156
6 8 19 0 0 8320 0 4 9 0 0 4
403 133
403 148
377 148
377 156
5 9 20 0 0 4224 0 4 9 0 0 4
397 133
397 148
386 148
386 156
4 10 21 0 0 4224 0 4 9 0 0 4
391 133
391 148
395 148
395 156
3 11 22 0 0 8320 0 4 9 0 0 4
385 133
385 148
404 148
404 156
2 12 23 0 0 8320 0 4 9 0 0 4
379 133
379 148
413 148
413 156
1 13 24 0 0 8320 0 4 9 0 0 4
373 133
373 148
422 148
422 156
7 7 25 0 0 8320 0 5 10 0 0 4
546 132
546 146
503 146
503 154
6 8 26 0 0 8320 0 5 10 0 0 4
540 132
540 146
512 146
512 154
5 9 27 0 0 4224 0 5 10 0 0 4
534 132
534 146
521 146
521 154
4 10 28 0 0 4224 0 5 10 0 0 4
528 132
528 146
530 146
530 154
3 11 29 0 0 8320 0 5 10 0 0 4
522 132
522 146
539 146
539 154
2 12 30 0 0 8320 0 5 10 0 0 4
516 132
516 146
548 146
548 154
1 13 31 0 0 8320 0 5 10 0 0 4
510 132
510 146
557 146
557 154
7 7 32 0 0 8320 0 6 11 0 0 4
679 135
679 145
638 145
638 153
6 8 33 0 0 8320 0 6 11 0 0 4
673 135
673 145
647 145
647 153
5 9 34 0 0 8320 0 6 11 0 0 4
667 135
667 145
656 145
656 153
4 10 35 0 0 4224 0 6 11 0 0 4
661 135
661 145
665 145
665 153
3 11 36 0 0 8320 0 6 11 0 0 4
655 135
655 145
674 145
674 153
2 12 37 0 0 8320 0 6 11 0 0 4
649 135
649 145
683 145
683 153
1 13 38 0 0 8320 0 6 11 0 0 4
643 135
643 145
692 145
692 153
7 7 39 0 0 8320 0 7 12 0 0 4
809 135
809 143
766 143
766 151
6 8 40 0 0 8320 0 7 12 0 0 4
803 135
803 143
775 143
775 151
5 9 41 0 0 8320 0 7 12 0 0 4
797 135
797 143
784 143
784 151
4 10 42 0 0 4224 0 7 12 0 0 4
791 135
791 143
793 143
793 151
3 11 43 0 0 8320 0 7 12 0 0 4
785 135
785 143
802 143
802 151
2 12 44 0 0 8320 0 7 12 0 0 4
779 135
779 143
811 143
811 151
1 13 45 0 0 8320 0 7 12 0 0 4
773 135
773 143
820 143
820 151
15 1 46 0 0 8320 0 30 8 0 0 3
283 346
221 346
221 223
16 2 47 0 0 8320 0 30 8 0 0 3
283 355
230 355
230 223
17 3 48 0 0 8320 0 30 8 0 0 3
283 364
239 364
239 223
18 4 49 0 0 8320 0 30 8 0 0 3
283 373
248 373
248 223
1 0 50 0 0 4224 0 9 0 0 76 2
368 226
368 346
2 0 51 0 0 4224 0 9 0 0 77 2
377 226
377 355
3 0 52 0 0 4224 0 9 0 0 78 2
386 226
386 364
4 0 53 0 0 4224 0 9 0 0 79 2
395 226
395 373
1 0 54 0 0 4224 0 10 0 0 80 2
503 224
503 348
2 0 55 0 0 4224 0 10 0 0 81 2
512 224
512 357
3 0 56 0 0 4224 0 10 0 0 82 2
521 224
521 366
4 0 57 0 0 4224 0 10 0 0 83 2
530 224
530 375
1 0 58 0 0 4224 0 11 0 0 84 2
638 223
638 349
2 0 59 0 0 4224 0 11 0 0 85 2
647 223
647 358
3 0 60 0 0 4224 0 11 0 0 86 2
656 223
656 367
4 0 61 0 0 4224 0 11 0 0 87 2
665 223
665 376
1 0 62 0 0 4224 0 12 0 0 88 4
766 221
766 335
768 335
768 350
2 0 63 0 0 4224 0 12 0 0 89 4
775 221
775 344
777 344
777 359
3 0 64 0 0 4224 0 12 0 0 90 4
784 221
784 353
786 353
786 368
4 0 65 0 0 4224 0 12 0 0 91 4
793 221
793 362
795 362
795 377
15 7 50 0 0 0 0 31 30 0 0 3
412 348
412 346
347 346
16 8 51 0 0 0 0 31 30 0 0 3
412 357
412 355
347 355
17 9 52 0 0 0 0 31 30 0 0 3
412 366
412 364
347 364
18 10 53 0 0 0 0 31 30 0 0 3
412 375
412 373
347 373
15 7 54 0 0 0 0 32 31 0 0 3
558 349
558 348
476 348
16 8 55 0 0 0 0 32 31 0 0 3
558 358
558 357
476 357
17 9 56 0 0 0 0 32 31 0 0 3
558 367
558 366
476 366
18 10 57 0 0 0 0 32 31 0 0 3
558 376
558 375
476 375
15 7 58 0 0 0 0 33 32 0 0 3
683 350
683 349
622 349
16 8 59 0 0 0 0 33 32 0 0 3
683 359
683 358
622 358
17 9 60 0 0 0 0 33 32 0 0 3
683 368
683 367
622 367
18 10 61 0 0 0 0 33 32 0 0 3
683 377
683 376
622 376
15 7 62 0 0 0 0 34 33 0 0 3
802 351
802 350
747 350
16 8 63 0 0 0 0 34 33 0 0 3
802 360
802 359
747 359
17 9 64 0 0 0 0 34 33 0 0 3
802 369
802 368
747 368
18 10 65 0 0 0 0 34 33 0 0 3
802 378
802 377
747 377
10 4 66 0 0 12416 0 34 23 0 0 5
866 378
949 378
949 430
760 430
760 454
3 3 67 0 0 4224 0 24 29 0 0 4
1164 501
1164 558
1173 558
1173 565
0 2 68 0 0 8192 0 0 29 121 0 3
1120 701
1182 701
1182 610
0 1 69 0 0 8192 0 0 29 107 0 4
936 770
936 668
1164 668
1164 610
4 3 70 0 0 8320 0 28 23 0 0 4
823 527
823 515
769 515
769 500
0 3 71 0 0 4096 0 0 28 105 0 3
710 633
832 633
832 579
0 2 72 0 0 4096 0 0 28 106 0 3
701 623
823 623
823 578
0 1 73 0 0 4096 0 0 28 111 0 3
888 606
814 606
814 579
2 4 74 0 0 4224 0 23 27 0 0 2
760 499
760 529
0 3 75 0 0 4224 0 0 27 132 0 3
991 750
769 750
769 581
0 2 72 0 0 0 0 0 27 106 0 3
701 612
760 612
760 580
0 1 69 0 0 0 0 0 27 107 0 3
692 605
751 605
751 581
1 4 76 0 0 8320 0 23 26 0 0 4
751 500
751 514
701 514
701 539
0 3 71 0 0 8192 0 0 26 109 0 3
908 790
710 790
710 584
0 2 72 0 0 4224 0 0 26 122 0 3
955 778
701 778
701 584
0 1 69 0 0 4224 0 0 26 129 0 3
937 770
692 770
692 584
1 4 77 0 0 4224 0 22 25 0 0 4
915 499
915 529
897 529
897 536
0 3 71 0 0 8320 0 0 25 131 0 3
973 790
906 790
906 581
2 2 78 0 0 8320 0 16 25 0 0 4
1074 721
1074 713
897 713
897 581
2 1 73 0 0 4224 0 15 25 0 0 3
1028 720
888 720
888 581
0 2 75 0 0 0 0 0 24 132 0 5
1025 671
1060 671
1060 550
1155 550
1155 500
0 1 79 0 0 4224 0 0 24 118 0 3
948 539
1146 539
1146 501
7 4 80 0 0 12416 0 34 24 0 0 5
866 351
976 351
976 438
1155 438
1155 455
3 9 81 0 0 16512 0 22 34 0 0 5
924 453
924 438
958 438
958 369
866 369
0 2 82 0 0 8192 0 0 22 117 0 5
967 451
953 451
953 506
933 506
933 499
8 3 82 0 0 8320 0 34 21 0 0 6
866 360
866 361
967 361
967 451
984 451
984 452
3 1 79 0 0 0 0 19 21 0 0 4
948 618
948 513
975 513
975 498
3 2 83 0 0 4224 0 20 21 0 0 4
1016 617
1016 509
993 509
993 498
0 1 69 0 0 0 0 0 20 129 0 2
1007 770
1007 662
2 2 68 0 0 8320 0 17 19 0 0 4
1120 723
1120 701
957 701
957 663
0 1 72 0 0 0 0 0 19 130 0 4
955 778
955 735
939 735
939 663
6 10 69 0 0 0 0 14 14 0 0 5
937 897
937 904
919 904
919 827
937 827
4 1 2 0 0 8320 0 14 18 0 0 4
964 891
964 902
984 902
984 908
1 3 2 0 0 0 0 18 14 0 0 4
984 908
984 903
973 903
973 891
1 2 2 0 0 0 0 18 14 0 0 4
984 908
984 903
982 903
982 891
1 1 2 0 0 0 0 18 14 0 0 4
984 908
984 903
991 903
991 891
3 5 3 0 0 0 0 13 14 0 0 3
1150 932
946 932
946 897
1 10 69 0 0 0 0 15 14 0 0 4
1028 756
1028 770
937 770
937 827
1 9 72 0 0 0 0 16 14 0 0 4
1074 757
1074 778
955 778
955 827
1 8 71 0 0 0 0 17 14 0 0 4
1120 759
1120 787
973 787
973 827
7 2 75 0 0 0 0 14 20 0 0 4
991 827
991 671
1025 671
1025 662
2
-27 0 0 0 700 0 0 0 0 3 2 1 34
5 Arial
0 0 0 25
1076 92 1348 177
1093 101 1352 165
25 SWARNENDU PAUL
19EE3FP18
-20 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 26
1094 176 1271 234
1108 185 1276 231
26 FP is shown as 00 
here.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
