CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 5 120 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
17
7 74LS165
97 421 392 0 14 29
0 8 8 34 35 36 37 2 2 3
5 2 4 38 3
0
0 0 13040 782
7 74LS165
-24 -60 25 -52
2 U1
54 -10 68 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 0 0 0
1 U
8953 0 0
0
0
9 Inverter~
13 320 328 0 2 22
0 9 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
4441 0 0
0
0
2 +V
167 892 472 0 1 3
0 18
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
9 2-In AND~
219 651 413 0 3 22
0 22 21 23
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6153 0 0
0
0
9 2-In NOR~
219 609 480 0 3 22
0 19 6 22
0
0 0 624 90
6 74LS02
-21 -24 21 -16
3 U7A
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5394 0 0
0
0
9 2-In AND~
219 687 476 0 3 22
0 7 20 21
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
9 CA 7-Seg~
184 892 93 0 18 19
10 10 11 12 13 14 15 16 39 17
0 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9914 0 0
0
0
10 Ascii Key~
169 420 278 0 11 12
0 37 36 35 34 40 41 42 9 0
0 56
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3747 0 0
0
0
7 74LS164
127 783 447 0 12 25
0 3 3 33 18 20 7 32 31 30
29 6 19
0
0 0 13040 90
7 74LS164
-24 -51 25 -43
2 U2
45 -6 59 2
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
7 Ground~
168 562 249 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
2 +V
167 517 244 0 1 3
0 8
0
0 0 54256 0
2 5V
6 -2 20 6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
7 Pulser~
4 175 532 0 10 12
0 43 44 4 45 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8903 0 0
0
0
7 Pulser~
4 903 416 0 10 12
0 46 47 33 48 0 0 5 5 5
7
0
0 0 4656 512
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3834 0 0
0
0
7 74LS273
150 774 322 0 18 37
0 24 23 49 50 32 31 30 29 51
52 53 54 28 27 26 25 55 56
0
0 0 13040 90
7 74LS273
-24 -60 25 -52
2 U4
54 -6 68 2
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
2 +V
167 689 59 0 1 3
0 24
0
0 0 54256 0
2 5V
-19 -2 -5 6
2 V4
-19 -12 -5 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
6 74LS47
187 804 242 0 14 29
0 28 27 26 25 57 58 16 15 14
13 12 11 10 59
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
9 Resistor~
219 750 36 0 3 5
0 24 17 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
42
2 0 3 0 0 4096 0 9 0 0 2 3
760 478
760 507
751 507
0 1 3 0 0 8320 0 0 9 4 0 4
462 446
462 529
751 529
751 478
11 1 2 0 0 12416 0 1 10 0 0 4
408 425
408 468
562 468
562 257
9 14 3 0 0 128 0 1 1 0 0 4
390 419
390 446
462 446
462 419
3 12 4 0 0 4224 0 12 1 0 0 3
199 523
417 523
417 419
2 10 5 0 0 4224 0 2 1 0 0 4
323 346
323 461
399 461
399 425
2 11 6 0 0 8320 0 5 9 0 0 6
624 499
624 586
848 586
848 383
805 383
805 414
6 1 7 0 0 12416 0 9 6 0 0 6
760 414
760 397
712 397
712 560
677 560
677 497
2 0 8 0 0 8192 0 1 0 0 21 4
408 355
408 333
517 333
517 325
7 0 2 0 0 128 0 1 0 0 3 3
453 355
453 345
562 345
8 1 9 0 0 4224 0 8 2 0 0 3
399 302
323 302
323 310
13 1 10 0 0 4224 0 16 7 0 0 4
823 209
823 152
871 152
871 129
12 2 11 0 0 8320 0 16 7 0 0 4
814 209
814 157
877 157
877 129
11 3 12 0 0 8320 0 16 7 0 0 4
805 209
805 162
883 162
883 129
10 4 13 0 0 8320 0 16 7 0 0 4
796 209
796 166
889 166
889 129
9 5 14 0 0 8320 0 16 7 0 0 4
787 209
787 174
895 174
895 129
8 6 15 0 0 8320 0 16 7 0 0 4
778 209
778 180
901 180
901 129
7 7 16 0 0 8320 0 7 16 0 0 4
907 129
907 185
769 185
769 209
2 9 17 0 0 4224 0 17 7 0 0 3
768 36
892 36
892 57
4 1 18 0 0 4224 0 9 3 0 0 3
796 484
892 484
892 481
1 1 8 0 0 8320 0 1 11 0 0 4
399 355
399 325
517 325
517 253
8 0 2 0 0 144 0 1 0 0 3 3
462 355
462 352
562 352
12 1 19 0 0 16512 0 9 5 0 0 6
814 414
814 396
836 396
836 573
606 573
606 499
5 2 20 0 0 12416 0 9 6 0 0 6
751 414
751 403
723 403
723 566
695 566
695 497
2 3 21 0 0 4224 0 4 6 0 0 3
659 434
686 434
686 452
1 3 22 0 0 4224 0 4 5 0 0 3
641 434
615 434
615 447
2 3 23 0 0 8320 0 14 4 0 0 3
742 353
742 389
650 389
1 0 24 0 0 8192 0 17 0 0 33 4
732 36
704 36
704 96
689 96
4 16 25 0 0 4224 0 16 14 0 0 2
796 279
796 289
3 15 26 0 0 4224 0 16 14 0 0 2
787 279
787 289
2 14 27 0 0 4224 0 16 14 0 0 2
778 279
778 289
1 13 28 0 0 4224 0 16 14 0 0 2
769 279
769 289
1 1 24 0 0 12416 0 14 15 0 0 4
733 359
733 363
689 363
689 68
8 10 29 0 0 4224 0 14 9 0 0 2
796 353
796 414
7 9 30 0 0 4224 0 14 9 0 0 2
787 353
787 414
6 8 31 0 0 4224 0 14 9 0 0 2
778 353
778 414
5 7 32 0 0 4224 0 14 9 0 0 2
769 353
769 414
3 3 33 0 0 8320 0 13 9 0 0 5
879 407
858 407
858 537
778 537
778 478
4 3 34 0 0 4224 0 8 1 0 0 4
423 302
423 349
417 349
417 355
3 4 35 0 0 4224 0 8 1 0 0 4
429 302
429 349
426 349
426 355
2 5 36 0 0 4224 0 8 1 0 0 2
435 302
435 355
1 6 37 0 0 8320 0 8 1 0 0 4
441 302
443 302
443 355
444 355
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
106 100 194 139
114 107 194 137
21 MODI OMKAR
19EE30018
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
