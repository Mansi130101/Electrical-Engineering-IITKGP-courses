CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 80 9
0 70 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1280 680
177209362 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 256 139 0 1 11
0 4
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
9 Inverter~
13 238 350 0 2 22
0 4 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7A
-30 2 -9 10
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
4441 0 0
0
0
14 Logic Display~
6 129 198 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
-24 2 -10 10
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 138 157 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 120 156 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
-24 2 -10 10
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
7 Ground~
168 96 89 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 396 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Pulser~
4 41 186 0 10 12
0 51 52 3 53 0 0 5 5 6
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3747 0 0
0
0
9 2-In AND~
219 414 109 0 3 22
0 6 30 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6D
8 16 29 24
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3549 0 0
0
0
9 2-In AND~
219 380 109 0 3 22
0 6 31 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6C
5 16 26 24
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
7931 0 0
0
0
9 2-In AND~
219 341 108 0 3 22
0 6 32 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6B
4 17 25 25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
9325 0 0
0
0
9 2-In AND~
219 305 109 0 3 22
0 6 33 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6A
5 16 26 24
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 383706678
65 0 0 0 4 1 1 0
1 U
8903 0 0
0
0
6 74LS47
187 409 638 0 14 29
0 23 24 25 36 54 55 43 41 42
40 39 38 37 56
0
0 0 13040 782
6 74LS47
-21 -60 21 -52
2 U2
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
9 CA 7-Seg~
184 291 641 0 18 19
10 37 38 39 40 42 41 43 57 35
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
28 30 63 38
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
9 CA 7-Seg~
184 68 640 0 18 19
10 44 45 46 47 49 48 50 58 35
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-62 -24 -27 -16
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7668 0 0
0
0
2 +V
167 68 514 0 1 3
0 34
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
6 74LS47
187 186 637 0 14 29
0 17 16 15 14 59 60 50 48 49
47 46 45 44 61
0
0 0 13040 782
6 74LS47
-21 -60 21 -52
2 U1
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
7 74LS273
150 282 412 0 18 37
0 5 3 18 19 20 21 22 23 24
25 17 16 15 14 23 24 25 36
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
6 74LS83
105 332 253 0 14 29
0 17 16 15 14 26 27 28 29 2
19 20 21 22 18
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
6 74LS95
110 157 105 0 12 25
0 4 3 3 13 12 11 10 2 6
7 8 9
0
0 0 13040 270
6 74LS95
-21 -51 21 -43
2 U3
45 0 59 8
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4871 0 0
0
0
8 Hex Key~
166 356 36 0 11 12
0 30 31 32 33 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3750 0 0
0
0
8 Hex Key~
166 144 42 0 11 12
0 13 12 11 10 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD1
-14 -37 14 -29
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8778 0 0
0
0
9 Resistor~
219 68 539 0 4 5
0 35 34 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
64
3 2 3 0 0 12416 0 8 18 0 0 5
65 177
94 177
94 277
250 277
250 385
1 1 4 0 0 8320 0 1 2 0 0 3
244 139
241 139
241 332
1 1 4 0 0 0 0 20 1 0 0 5
183 78
183 68
241 68
241 139
244 139
2 1 5 0 0 4224 0 2 18 0 0 2
241 368
241 379
9 0 6 0 0 12416 0 20 0 0 35 4
147 142
227 142
227 78
312 78
1 10 7 0 0 12416 0 4 20 0 0 4
138 143
138 150
138 150
138 142
1 11 8 0 0 4224 0 3 20 0 0 2
129 184
129 142
1 12 9 0 0 0 0 5 20 0 0 2
120 142
120 142
1 8 2 0 0 8320 0 6 20 0 0 4
96 83
96 64
120 64
120 78
7 4 10 0 0 4224 0 20 22 0 0 5
129 78
129 66
137 66
137 66
135 66
6 3 11 0 0 12416 0 20 22 0 0 4
138 78
138 74
141 74
141 66
5 2 12 0 0 4224 0 20 22 0 0 2
147 78
147 66
4 1 13 0 0 4224 0 20 22 0 0 3
156 78
156 66
153 66
2 0 3 0 0 0 0 20 0 0 15 2
174 72
174 64
3 3 3 0 0 0 0 8 20 0 0 5
65 177
203 177
203 64
165 64
165 72
9 1 2 0 0 0 0 19 7 0 0 4
375 223
375 222
396 222
396 224
1 0 6 0 0 0 0 9 0 0 34 3
421 87
421 78
387 78
0 4 14 0 0 8320 0 0 19 42 0 5
286 501
159 501
159 192
321 192
321 223
0 3 15 0 0 8320 0 0 19 43 0 5
277 490
171 490
171 203
312 203
312 223
0 2 16 0 0 8320 0 0 19 44 0 5
268 477
182 477
182 213
303 213
303 223
0 1 17 0 0 8320 0 0 19 45 0 4
259 462
192 462
192 223
294 223
14 3 18 0 0 8320 0 19 18 0 0 4
375 287
375 300
259 300
259 385
10 4 19 0 0 12416 0 19 18 0 0 4
321 287
321 308
268 308
268 385
11 5 20 0 0 12416 0 19 18 0 0 4
330 287
330 317
277 317
277 385
12 6 21 0 0 12416 0 19 18 0 0 4
339 287
339 328
286 328
286 385
13 7 22 0 0 12416 0 19 18 0 0 5
348 287
347 287
347 337
295 337
295 385
0 8 23 0 0 8192 0 0 18 46 0 5
295 487
355 487
355 351
304 351
304 385
0 9 24 0 0 8192 0 0 18 47 0 5
304 476
346 476
346 361
313 361
313 385
0 10 25 0 0 8192 0 0 18 48 0 5
313 462
337 462
337 371
322 371
322 385
3 5 26 0 0 12416 0 12 19 0 0 4
303 132
303 147
330 147
330 223
3 6 27 0 0 4224 0 11 19 0 0 2
339 131
339 223
3 7 28 0 0 4224 0 10 19 0 0 4
378 132
378 201
348 201
348 223
3 8 29 0 0 4224 0 9 19 0 0 4
412 132
412 212
357 212
357 223
0 1 6 0 0 0 0 0 10 35 0 3
349 78
387 78
387 87
1 1 6 0 0 0 0 12 11 0 0 6
312 87
312 78
349 78
349 78
348 78
348 86
2 1 30 0 0 8320 0 9 21 0 0 3
403 87
403 60
365 60
2 2 31 0 0 4224 0 10 21 0 0 4
369 87
369 68
359 68
359 60
2 3 32 0 0 8320 0 11 21 0 0 4
330 86
330 68
353 68
353 60
2 4 33 0 0 8320 0 12 21 0 0 4
294 87
294 59
347 59
347 60
2 1 34 0 0 4224 0 23 16 0 0 2
68 521
68 523
9 9 35 0 0 8320 0 14 15 0 0 4
291 605
291 580
68 580
68 604
14 4 14 0 0 0 0 18 17 0 0 4
286 449
286 594
178 594
178 604
13 3 15 0 0 0 0 18 17 0 0 4
277 449
277 586
169 586
169 604
12 2 16 0 0 0 0 18 17 0 0 4
268 449
268 572
160 572
160 604
11 1 17 0 0 0 0 18 17 0 0 4
259 449
259 566
151 566
151 604
15 1 23 0 0 4224 0 18 13 0 0 4
295 449
295 586
374 586
374 605
16 2 24 0 0 4224 0 18 13 0 0 4
304 449
304 580
383 580
383 605
17 3 25 0 0 4224 0 18 13 0 0 4
313 449
313 574
392 574
392 605
18 4 36 0 0 4224 0 18 13 0 0 4
322 449
322 568
401 568
401 605
1 13 37 0 0 8320 0 14 13 0 0 4
270 677
270 686
428 686
428 675
12 2 38 0 0 8320 0 13 14 0 0 4
419 675
419 685
276 685
276 677
11 3 39 0 0 8320 0 13 14 0 0 4
410 675
410 685
282 685
282 677
10 4 40 0 0 8320 0 13 14 0 0 4
401 675
401 685
288 685
288 677
8 6 41 0 0 8320 0 13 14 0 0 4
383 675
383 685
300 685
300 677
9 5 42 0 0 8320 0 13 14 0 0 4
392 675
392 685
294 685
294 677
7 7 43 0 0 8320 0 13 14 0 0 4
374 675
374 685
306 685
306 677
1 13 44 0 0 8320 0 15 17 0 0 4
47 676
47 685
205 685
205 674
12 2 45 0 0 8320 0 17 15 0 0 4
196 674
196 684
53 684
53 676
11 3 46 0 0 8320 0 17 15 0 0 4
187 674
187 684
59 684
59 676
10 4 47 0 0 8320 0 17 15 0 0 4
178 674
178 684
65 684
65 676
8 6 48 0 0 8320 0 17 15 0 0 4
160 674
160 684
77 684
77 676
9 5 49 0 0 8320 0 17 15 0 0 4
169 674
169 684
71 684
71 676
7 7 50 0 0 8320 0 17 15 0 0 4
151 674
151 684
83 684
83 676
1 9 35 0 0 0 0 23 15 0 0 2
68 557
68 604
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 74
481 187 699 267
491 197 701 257
74 4-bit multiplier; using the 
shifter and adder to multiply 
the digits
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
