CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
390 140 20 200 9
48 116 1872 995
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 116 1872 995
143654930 0
0
6 Title:
5 Name:
0
0
0
19
9 2-In AND~
219 851 349 0 3 22
0 29 28 4
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U5C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
8953 0 0
0
0
9 2-In NOR~
219 927 351 0 3 22
0 30 31 5
0
0 0 624 90
6 74LS02
-21 -24 21 -16
3 U4A
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
4441 0 0
0
0
7 Ground~
168 729 372 0 1 3
0 2
0
0 0 53360 782
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 616 366 0 1 3
0 33
0
0 0 54256 782
2 5V
-8 -15 6 -7
2 V3
-8 -25 6 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
2 +V
167 964 200 0 1 3
0 7
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
9 Inverter~
13 573 380 0 2 22
0 10 8
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
-31 -11 -10 -3
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
7734 0 0
0
0
2 +V
167 1064 173 0 1 3
0 3
0
0 0 54256 90
2 5V
-7 -15 7 -7
2 V6
-7 -25 7 -17
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
6 74LS47
187 1084 313 0 14 29
0 19 20 21 22 53 54 12 13 14
15 16 17 18 55
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
9 CA 7-Seg~
184 1155 232 0 18 19
10 18 17 16 15 14 13 12 56 11
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
7 74LS165
97 664 420 0 14 29
0 33 33 34 35 36 37 2 2 6
8 2 38 57 6
0
0 0 13040 782
7 74LS165
-24 -60 25 -52
2 U7
54 -10 68 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 74LS273
150 1007 259 0 18 37
0 7 27 58 59 60 61 23 24 25
26 62 63 64 65 19 20 21 22
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
7 74LS164
127 899 415 0 12 25
0 6 6 32 9 29 28 23 24 25
26 30 31
0
0 0 13040 90
7 74LS164
-24 -51 25 -43
2 U1
45 -6 59 2
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
7 Ground~
168 641 486 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3834 0 0
0
0
7 Pulser~
4 507 478 0 10 12
0 66 67 38 68 0 0 20 20 21
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3363 0 0
0
0
10 Ascii Key~
169 662 284 0 11 12
0 37 36 35 34 69 70 71 10 0
0 56
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
7668 0 0
0
0
7 Pulser~
4 1038 476 0 10 12
0 72 73 32 74 0 0 20 20 21
7
0
0 0 4656 512
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4718 0 0
0
0
2 +V
167 913 495 0 1 3
0 9
0
0 0 54256 180
2 5V
7 -2 21 6
2 V5
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3874 0 0
0
0
9 2-In AND~
219 894 224 0 3 22
0 4 5 27
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U5B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
6671 0 0
0
0
9 Resistor~
219 1115 171 0 3 5
0 3 11 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
42
3 1 4 0 0 4224 0 1 18 0 0 3
850 325
850 245
884 245
3 2 5 0 0 4224 0 2 18 0 0 3
933 318
933 245
902 245
9 0 6 0 0 8192 0 10 0 0 9 3
633 447
633 515
705 515
8 0 2 0 0 4096 0 10 0 0 5 2
705 383
705 373
1 7 2 0 0 4096 0 3 10 0 0 3
722 373
696 373
696 383
1 1 7 0 0 8320 0 11 5 0 0 3
969 223
964 223
964 209
11 1 2 0 0 4224 0 10 13 0 0 3
651 453
651 480
641 480
10 2 8 0 0 8320 0 10 6 0 0 4
642 453
642 460
576 460
576 398
14 1 6 0 0 8320 0 10 12 0 0 4
705 447
705 515
867 515
867 446
4 1 9 0 0 8320 0 12 17 0 0 3
912 452
913 452
913 480
8 1 10 0 0 4224 0 15 6 0 0 3
641 308
576 308
576 362
1 1 3 0 0 4224 0 19 7 0 0 2
1097 171
1075 171
2 9 11 0 0 8320 0 19 9 0 0 3
1133 171
1155 171
1155 196
7 7 12 0 0 4224 0 8 9 0 0 3
1122 277
1170 277
1170 268
8 6 13 0 0 4224 0 8 9 0 0 3
1122 286
1164 286
1164 268
9 5 14 0 0 4224 0 8 9 0 0 3
1122 295
1158 295
1158 268
10 4 15 0 0 8320 0 8 9 0 0 3
1122 304
1152 304
1152 268
11 3 16 0 0 8320 0 8 9 0 0 3
1122 313
1146 313
1146 268
12 2 17 0 0 8320 0 8 9 0 0 3
1122 322
1140 322
1140 268
13 1 18 0 0 8320 0 8 9 0 0 3
1122 331
1134 331
1134 268
1 15 19 0 0 4224 0 8 11 0 0 2
1052 277
1039 277
2 16 20 0 0 4224 0 8 11 0 0 2
1052 286
1039 286
3 17 21 0 0 4224 0 8 11 0 0 2
1052 295
1039 295
4 18 22 0 0 4224 0 8 11 0 0 2
1052 304
1039 304
7 7 23 0 0 4224 0 12 11 0 0 3
885 382
885 277
975 277
8 8 24 0 0 4224 0 12 11 0 0 3
894 382
894 286
975 286
9 9 25 0 0 4224 0 12 11 0 0 3
903 382
903 295
975 295
10 10 26 0 0 4224 0 12 11 0 0 3
912 382
912 304
975 304
3 2 27 0 0 4224 0 18 11 0 0 4
893 200
952 200
952 232
975 232
6 2 28 0 0 8320 0 12 1 0 0 4
876 382
876 371
859 371
859 370
5 1 29 0 0 4224 0 12 1 0 0 3
867 382
841 382
841 370
1 11 30 0 0 4224 0 2 12 0 0 3
924 370
924 382
921 382
2 12 31 0 0 4224 0 2 12 0 0 3
942 370
942 382
930 382
3 3 32 0 0 4224 0 16 12 0 0 3
1014 467
894 467
894 446
1 0 33 0 0 4096 0 10 0 0 36 2
642 383
642 365
2 1 33 0 0 16512 0 10 4 0 0 5
651 383
651 382
650 382
650 365
626 365
2 0 6 0 0 0 0 12 0 0 9 3
876 446
876 461
867 461
4 3 34 0 0 4224 0 15 10 0 0 4
665 308
665 374
660 374
660 383
3 4 35 0 0 4224 0 15 10 0 0 4
671 308
671 374
669 374
669 383
2 5 36 0 0 4224 0 15 10 0 0 4
677 308
677 374
678 374
678 383
1 6 37 0 0 4224 0 15 10 0 0 4
683 308
683 374
687 374
687 383
12 3 38 0 0 8320 0 10 14 0 0 3
660 447
660 469
531 469
1
-20 0 0 0 400 0 0 0 0 3 2 1 34
6 Gadugi
0 0 0 25
668 179 855 242
674 184 848 232
25 SWARNENDU PAUL
19EE3FP18
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
