CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 330 1 100 9
0 80 1544 832
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 80 1544 832
143654930 0
0
6 Title:
5 Name:
0
0
0
45
7 Ground~
168 375 570 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 74LS173
129 305 548 0 14 29
0 2 2 2 3 17 16 15 14 2
2 10 11 12 13
0
0 0 13024 602
7 74LS173
-24 -51 25 -43
3 U19
47 -3 68 5
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4441 0 0
0
0
9 CA 7-Seg~
184 284 381 0 18 19
10 24 23 22 21 20 19 18 85 9
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3618 0 0
0
0
6 74LS47
187 270 459 0 14 29
0 10 11 12 13 86 87 18 19 20
21 22 23 24 88
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
3 U14
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
6 74LS47
187 454 511 0 14 29
0 17 16 15 14 89 90 25 26 27
28 29 30 31 91
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
3 U13
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
9 CA 7-Seg~
184 468 433 0 18 19
10 31 30 29 28 27 26 25 92 8
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7734 0 0
0
0
7 Ground~
168 590 642 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 74LS173
129 502 611 0 14 29
0 2 2 2 3 35 34 33 32 2
2 17 16 15 14
0
0 0 13024 602
7 74LS173
-24 -51 25 -43
3 U18
47 -3 68 5
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
9 CA 7-Seg~
184 648 476 0 18 19
10 42 41 40 39 38 37 36 93 7
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3549 0 0
0
0
6 74LS47
187 634 554 0 14 29
0 35 34 33 32 94 95 36 37 38
39 40 41 42 96
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
3 U17
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 Ground~
168 747 660 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 933 669 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 74LS173
129 682 647 0 14 29
0 2 2 2 3 45 45 44 43 2
2 35 34 33 32
0
0 0 13024 602
7 74LS173
-24 -51 25 -43
3 U15
47 -3 68 5
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
2 +V
167 987 243 0 1 3
0 4
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
2 +V
167 731 823 0 1 3
0 77
0
0 0 54240 180
2 5V
7 -2 21 6
2 V3
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Pulser~
4 817 1267 0 10 12
0 97 98 76 3 0 0 7 7 8
7
0
0 0 4640 90
0
2 V1
23 -5 37 3
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
6 74LS47
187 1013 758 0 14 29
0 47 48 49 50 77 76 78 79 80
81 82 83 84 76
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
9 CA 7-Seg~
184 1008 529 0 18 19
10 84 83 82 81 80 79 78 99 5
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6671 0 0
0
0
6 74LS93
109 818 1165 0 8 17
0 60 59 76 58 60 68 59 58
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
5 4073~
219 692 938 0 4 22
0 59 61 64 67
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U9B
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 7 0
1 U
4871 0 0
0
0
8 2-In OR~
219 572 880 0 3 22
0 72 71 50
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U10B
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 8 0
1 U
3750 0 0
0
0
8 3-In OR~
219 1145 893 0 4 22
0 75 74 73 47
0
0 0 608 90
4 4075
-14 -24 14 -16
3 U5A
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 3 0
1 U
8778 0 0
0
0
9 Inverter~
13 872 1050 0 2 22
0 60 64
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
538 0 0
0
0
9 Inverter~
13 755 1052 0 2 22
0 58 63
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U3D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
6843 0 0
0
0
9 Inverter~
13 793 1051 0 2 22
0 59 62
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U3C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3136 0 0
0
0
9 Inverter~
13 832 1051 0 2 22
0 68 61
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U3B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
5950 0 0
0
0
5 4073~
219 1063 968 0 4 22
0 60 62 61 75
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U9C
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 7 0
1 U
5670 0 0
0
0
5 4073~
219 1155 967 0 4 22
0 59 64 61 74
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U4A
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 9 0
1 U
6828 0 0
0
0
5 4073~
219 1247 967 0 4 22
0 58 61 64 73
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U4B
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 9 0
1 U
6735 0 0
0
0
5 4073~
219 911 940 0 4 22
0 59 61 64 70
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U4C
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 9 0
1 U
8365 0 0
0
0
9 4-In AND~
219 974 937 0 5 22
0 58 60 62 61 69
0
0 0 608 90
6 74LS21
-21 -28 21 -20
3 U8A
19 -5 40 3
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 1 10 0
1 U
4132 0 0
0
0
8 2-In OR~
219 934 880 0 3 22
0 70 69 48
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U10C
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 8 0
1 U
4551 0 0
0
0
9 4-In AND~
219 752 936 0 5 22
0 63 62 68 64 66
0
0 0 608 90
6 74LS21
-21 -28 21 -20
3 U8B
19 -5 40 3
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 2 10 0
1 U
3635 0 0
0
0
9 4-In AND~
219 817 935 0 5 22
0 58 62 61 60 65
0
0 0 608 90
6 74LS21
-21 -28 21 -20
3 U7A
19 -5 40 3
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 1 5 0
1 U
3973 0 0
0
0
8 3-In OR~
219 730 880 0 4 22
0 67 66 65 49
0
0 0 608 90
4 4075
-14 -24 14 -16
3 U5B
28 -3 49 5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 3 0
1 U
3851 0 0
0
0
5 4073~
219 530 949 0 4 22
0 58 61 62 72
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U6A
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
8383 0 0
0
0
5 4073~
219 593 956 0 4 22
0 63 62 64 71
0
0 0 608 90
4 4073
-7 -24 21 -16
4 U11A
13 -5 41 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 11 0
1 U
9334 0 0
0
0
9 CA 7-Seg~
184 830 527 0 18 19
10 57 56 55 54 53 52 51 100 6
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7471 0 0
0
0
6 74LS47
187 816 605 0 14 29
0 45 46 44 43 101 102 51 52 53
54 55 56 57 103
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
3 U12
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3334 0 0
0
0
7 74LS173
129 868 708 0 14 29
0 2 2 2 3 47 48 49 50 2
2 45 46 44 43
0
0 0 13024 602
7 74LS173
-24 -51 25 -43
3 U16
47 -3 68 5
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3559 0 0
0
0
9 Resistor~
219 284 316 0 4 5
0 9 4 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 469 370 0 4 5
0 8 4 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 648 410 0 4 5
0 7 4 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 830 456 0 4 5
0 6 4 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 987 432 0 4 5
0 5 4 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7939 0 0
0
0
159
0 4 3 0 0 4096 0 0 2 4 0 4
324 739
324 596
307 596
307 582
0 4 3 0 0 0 0 0 8 4 0 2
504 739
504 645
0 4 3 0 0 8192 0 0 40 4 0 4
683 739
683 756
870 756
870 742
4 4 3 0 0 8336 0 16 13 0 0 6
817 1237
817 1205
320 1205
320 739
684 739
684 681
2 0 4 0 0 4096 0 44 0 0 8 2
830 438
830 294
2 0 4 0 0 0 0 43 0 0 8 2
648 392
648 294
2 0 4 0 0 0 0 42 0 0 8 2
469 352
469 294
2 0 4 0 0 8320 0 41 0 0 9 3
284 298
284 294
987 294
1 2 4 0 0 0 0 14 45 0 0 2
987 252
987 414
1 9 5 0 0 4224 0 45 18 0 0 4
987 450
987 485
1008 485
1008 493
1 9 6 0 0 4224 0 44 38 0 0 2
830 474
830 491
1 9 7 0 0 4224 0 43 9 0 0 2
648 428
648 440
1 9 8 0 0 4224 0 42 6 0 0 3
469 388
469 397
468 397
1 9 9 0 0 4224 0 41 3 0 0 2
284 334
284 345
3 2 2 0 0 4096 0 2 2 0 0 2
316 588
325 588
2 0 2 0 0 0 0 2 0 0 17 3
325 588
325 589
334 589
1 0 2 0 0 12288 0 2 0 0 19 5
334 582
334 592
361 592
361 557
375 557
10 0 2 0 0 0 0 2 0 0 19 3
325 512
325 508
334 508
9 1 2 0 0 12288 0 2 1 0 0 4
334 512
334 508
375 508
375 564
11 1 10 0 0 4224 0 2 4 0 0 4
298 518
298 504
311 504
311 496
12 2 11 0 0 4224 0 2 4 0 0 4
289 518
289 504
302 504
302 496
13 3 12 0 0 4224 0 2 4 0 0 4
280 518
280 504
293 504
293 496
14 4 13 0 0 4224 0 2 4 0 0 4
271 518
271 504
284 504
284 496
0 8 14 0 0 12416 0 0 2 31 0 5
468 553
435 553
435 655
271 655
271 582
0 7 15 0 0 12416 0 0 2 30 0 5
477 558
422 558
422 645
280 645
280 582
0 6 16 0 0 12416 0 0 2 29 0 5
486 569
408 569
408 640
289 640
289 582
0 5 17 0 0 20608 0 0 2 28 0 7
495 576
429 576
429 577
399 577
399 634
298 634
298 582
11 1 17 0 0 0 0 8 5 0 0 2
495 581
495 548
12 2 16 0 0 0 0 8 5 0 0 2
486 581
486 548
13 3 15 0 0 0 0 8 5 0 0 2
477 581
477 548
14 4 14 0 0 0 0 8 5 0 0 2
468 581
468 548
7 7 18 0 0 8320 0 4 3 0 0 3
311 426
311 417
299 417
8 6 19 0 0 4224 0 4 3 0 0 3
302 426
302 417
293 417
9 5 20 0 0 4224 0 4 3 0 0 3
293 426
293 417
287 417
10 4 21 0 0 4224 0 4 3 0 0 3
284 426
284 417
281 417
11 3 22 0 0 4224 0 4 3 0 0 2
275 426
275 417
12 2 23 0 0 4224 0 4 3 0 0 4
266 426
266 420
269 420
269 417
13 1 24 0 0 4224 0 4 3 0 0 3
257 426
257 417
263 417
7 7 25 0 0 8320 0 5 6 0 0 3
495 478
495 469
483 469
8 6 26 0 0 4224 0 5 6 0 0 3
486 478
486 469
477 469
9 5 27 0 0 4224 0 5 6 0 0 3
477 478
477 469
471 469
10 4 28 0 0 4224 0 5 6 0 0 3
468 478
468 469
465 469
11 3 29 0 0 4224 0 5 6 0 0 2
459 478
459 469
12 2 30 0 0 4224 0 5 6 0 0 4
450 478
450 472
453 472
453 469
13 1 31 0 0 4224 0 5 6 0 0 3
441 478
441 469
447 469
3 2 2 0 0 0 0 8 8 0 0 2
513 651
522 651
2 0 2 0 0 0 0 8 0 0 48 2
522 651
531 651
1 0 2 0 0 0 0 8 0 0 50 5
531 645
531 654
576 654
576 627
590 627
10 0 2 0 0 0 0 8 0 0 50 3
522 575
522 571
536 571
9 1 2 0 0 0 0 8 7 0 0 6
531 575
531 571
580 571
580 596
590 596
590 636
0 8 32 0 0 4224 0 0 8 65 0 5
648 598
550 598
550 659
468 659
468 645
0 7 33 0 0 4224 0 0 8 64 0 5
657 603
550 603
550 659
477 659
477 645
0 6 34 0 0 12416 0 0 8 63 0 5
667 609
611 609
611 709
486 709
486 645
0 5 35 0 0 12416 0 0 8 62 0 5
676 611
617 611
617 703
495 703
495 645
7 7 36 0 0 8320 0 10 9 0 0 3
675 521
675 512
663 512
8 6 37 0 0 4224 0 10 9 0 0 3
666 521
666 512
657 512
9 5 38 0 0 4224 0 10 9 0 0 3
657 521
657 512
651 512
10 4 39 0 0 4224 0 10 9 0 0 3
648 521
648 512
645 512
11 3 40 0 0 4224 0 10 9 0 0 2
639 521
639 512
12 2 41 0 0 4224 0 10 9 0 0 4
630 521
630 515
633 515
633 512
13 1 42 0 0 4224 0 10 9 0 0 3
621 521
621 512
627 512
11 1 35 0 0 0 0 13 10 0 0 5
675 617
676 617
676 609
675 609
675 591
12 2 34 0 0 0 0 13 10 0 0 5
666 617
667 617
667 609
666 609
666 591
13 3 33 0 0 0 0 13 10 0 0 5
657 617
658 617
658 609
657 609
657 591
14 4 32 0 0 0 0 13 10 0 0 5
648 617
649 617
649 609
648 609
648 591
0 8 43 0 0 12416 0 0 13 83 0 5
834 658
760 658
760 695
648 695
648 681
0 7 44 0 0 12416 0 0 13 82 0 5
843 662
760 662
760 695
657 695
657 681
0 6 45 0 0 16384 0 0 13 69 0 6
853 675
853 668
760 668
760 692
666 692
666 681
0 5 45 0 0 4224 0 0 13 80 0 5
861 675
760 675
760 695
675 695
675 681
3 0 2 0 0 0 0 13 0 0 71 3
693 687
693 691
702 691
2 0 2 0 0 0 0 13 0 0 74 3
702 687
702 691
711 691
10 0 2 0 0 0 0 13 0 0 73 3
702 611
702 607
711 607
9 0 2 0 0 0 0 13 0 0 74 4
711 611
711 607
747 607
747 646
1 1 2 0 0 0 0 13 11 0 0 6
711 681
711 691
733 691
733 646
747 646
747 654
3 0 2 0 0 0 0 40 0 0 76 3
879 748
879 752
891 752
2 0 2 0 0 0 0 40 0 0 77 3
888 748
888 752
901 752
1 0 2 0 0 12416 0 40 0 0 78 4
897 742
897 752
917 752
917 655
9 1 2 0 0 0 0 40 12 0 0 4
897 672
897 655
933 655
933 663
10 1 2 0 0 0 0 40 12 0 0 4
888 672
888 655
933 655
933 663
11 1 45 0 0 0 0 40 39 0 0 4
861 678
861 650
857 650
857 642
12 2 46 0 0 4224 0 40 39 0 0 4
852 678
852 650
848 650
848 642
13 3 44 0 0 0 0 40 39 0 0 4
843 678
843 650
839 650
839 642
14 4 43 0 0 0 0 40 39 0 0 4
834 678
834 650
830 650
830 642
0 5 47 0 0 8320 0 0 40 145 0 4
1065 807
1065 799
861 799
861 742
0 6 48 0 0 8192 0 0 40 128 0 4
937 833
937 771
852 771
852 742
0 7 49 0 0 4096 0 0 40 118 0 4
843 840
843 740
843 740
843 742
0 8 50 0 0 12288 0 0 40 142 0 4
833 818
833 803
834 803
834 742
7 7 51 0 0 8320 0 39 38 0 0 3
857 572
857 563
845 563
8 6 52 0 0 4224 0 39 38 0 0 3
848 572
848 563
839 563
9 5 53 0 0 4224 0 39 38 0 0 3
839 572
839 563
833 563
10 4 54 0 0 4224 0 39 38 0 0 3
830 572
830 563
827 563
11 3 55 0 0 4224 0 39 38 0 0 2
821 572
821 563
12 2 56 0 0 4224 0 39 38 0 0 4
812 572
812 566
815 566
815 563
13 1 57 0 0 4224 0 39 38 0 0 3
803 572
803 563
809 563
4 0 58 0 0 12288 0 19 0 0 98 4
798 1201
798 1205
771 1205
771 1111
2 0 59 0 0 12288 0 19 0 0 139 5
816 1195
816 1212
783 1212
783 1126
807 1126
1 0 60 0 0 12288 0 19 0 0 141 5
825 1195
825 1205
847 1205
847 1117
825 1117
0 1 58 0 0 4096 0 0 36 138 0 3
798 1111
520 1111
520 970
0 2 61 0 0 4096 0 0 36 109 0 3
821 1003
529 1003
529 970
0 3 62 0 0 4096 0 0 36 102 0 3
593 1023
538 1023
538 970
0 1 63 0 0 4224 0 0 37 111 0 3
738 995
583 995
583 977
0 2 62 0 0 4096 0 0 37 112 0 3
750 1023
592 1023
592 977
0 3 64 0 0 8192 0 0 37 114 0 4
766 994
766 1013
601 1013
601 977
5 3 65 0 0 8320 0 34 35 0 0 4
816 911
816 903
742 903
742 896
5 2 66 0 0 12416 0 33 35 0 0 4
751 912
751 925
733 925
733 895
4 1 67 0 0 8320 0 20 35 0 0 4
691 914
691 911
724 911
724 896
0 1 58 0 0 0 0 0 34 138 0 6
771 1078
771 1073
772 1073
772 967
803 967
803 956
0 2 62 0 0 0 0 0 34 130 0 2
812 1013
812 956
0 3 61 0 0 0 0 0 34 136 0 3
835 1023
821 1023
821 956
0 4 60 0 0 4096 0 0 34 141 0 4
858 1095
858 965
830 965
830 956
2 1 63 0 0 0 0 24 33 0 0 3
758 1034
738 1034
738 957
0 2 62 0 0 0 0 0 33 130 0 4
796 1023
749 1023
749 957
747 957
0 3 68 0 0 8320 0 0 33 140 0 5
816 1093
743 1093
743 964
756 964
756 957
0 4 64 0 0 0 0 0 33 117 0 3
892 994
765 994
765 957
0 1 59 0 0 8192 0 0 20 139 0 3
807 1099
682 1099
682 959
0 2 61 0 0 0 0 0 20 136 0 4
887 1020
887 984
691 984
691 959
0 3 64 0 0 8192 0 0 20 137 0 4
892 1030
892 975
700 975
700 959
3 4 49 0 0 8320 0 17 35 0 0 4
1036 795
1036 840
733 840
733 850
5 2 69 0 0 8320 0 31 32 0 0 4
973 913
973 909
946 909
946 896
4 1 70 0 0 8320 0 30 32 0 0 4
910 916
910 911
928 911
928 896
0 1 59 0 0 4096 0 0 30 132 0 2
901 1111
901 961
0 2 61 0 0 0 0 0 30 136 0 2
910 1020
910 961
0 3 64 0 0 0 0 0 30 137 0 2
919 1030
919 961
0 1 58 0 0 0 0 0 31 135 0 2
960 1121
960 958
0 2 60 0 0 4096 0 0 31 129 0 2
969 1105
969 958
0 3 62 0 0 0 0 0 31 130 0 2
978 1013
978 958
0 4 61 0 0 0 0 0 31 136 0 2
987 1020
987 958
2 3 48 0 0 8320 0 17 32 0 0 4
1045 795
1045 833
937 833
937 850
0 1 60 0 0 4224 0 0 27 141 0 3
825 1105
1053 1105
1053 989
2 2 62 0 0 8320 0 25 27 0 0 4
796 1033
796 1013
1062 1013
1062 989
0 3 61 0 0 0 0 0 27 136 0 2
1071 1020
1071 989
0 1 59 0 0 4224 0 0 28 139 0 3
807 1111
1145 1111
1145 988
0 2 64 0 0 0 0 0 28 137 0 2
1154 1030
1154 988
0 3 61 0 0 0 0 0 28 136 0 2
1163 1020
1163 988
0 1 58 0 0 4224 0 0 29 138 0 3
798 1121
1237 1121
1237 988
2 2 61 0 0 8320 0 26 29 0 0 4
835 1033
835 1020
1246 1020
1246 988
2 3 64 0 0 8320 0 23 29 0 0 4
875 1032
875 1030
1255 1030
1255 988
8 1 58 0 0 0 0 19 24 0 0 4
798 1131
798 1078
758 1078
758 1070
7 1 59 0 0 0 0 19 25 0 0 4
807 1131
807 1075
796 1075
796 1069
6 1 68 0 0 0 0 19 26 0 0 4
816 1131
816 1084
835 1084
835 1069
5 1 60 0 0 0 0 19 23 0 0 4
825 1131
825 1095
875 1095
875 1068
3 4 50 0 0 8320 0 21 17 0 0 4
575 850
575 818
1027 818
1027 795
4 2 71 0 0 12416 0 37 21 0 0 4
592 932
592 919
584 919
584 896
4 1 72 0 0 8320 0 36 21 0 0 4
529 925
529 919
566 919
566 896
4 1 47 0 0 0 0 22 17 0 0 4
1148 863
1148 807
1054 807
1054 795
4 3 73 0 0 8320 0 29 22 0 0 4
1246 943
1246 924
1157 924
1157 909
4 2 74 0 0 4224 0 28 22 0 0 4
1154 943
1154 924
1148 924
1148 908
4 1 75 0 0 8320 0 27 22 0 0 4
1062 944
1062 924
1139 924
1139 909
14 0 76 0 0 12288 0 17 0 0 150 5
973 731
943 731
943 782
689 782
689 801
6 3 76 0 0 16512 0 17 16 0 0 8
973 795
689 795
689 801
508 801
508 1259
781 1259
781 1243
808 1243
1 5 77 0 0 8320 0 15 17 0 0 3
731 808
731 795
982 795
7 7 78 0 0 4224 0 18 17 0 0 4
1023 565
1023 706
1054 706
1054 725
8 6 79 0 0 12416 0 17 18 0 0 4
1045 725
1045 710
1017 710
1017 565
9 5 80 0 0 12416 0 17 18 0 0 4
1036 725
1036 715
1011 715
1011 565
10 4 81 0 0 12416 0 17 18 0 0 4
1027 725
1027 720
1005 720
1005 565
11 3 82 0 0 8320 0 17 18 0 0 3
1018 725
999 725
999 565
12 2 83 0 0 8320 0 17 18 0 0 4
1009 725
994 725
994 565
993 565
13 1 84 0 0 12416 0 17 18 0 0 4
1000 725
1000 710
987 710
987 565
3 3 76 0 0 0 0 16 19 0 0 4
808 1243
808 1203
807 1203
807 1201
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
