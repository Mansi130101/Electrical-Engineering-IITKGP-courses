CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
3 86 1283 695
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
3 86 1283 695
143654930 0
0
6 Title:
5 Name:
0
0
0
9
14 Logic Display~
6 431 285 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
7 Ground~
168 351 237 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
9 CA 7-Seg~
184 555 105 0 18 19
10 9 8 7 6 5 10 11 25 4
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3618 0 0
0
0
2 +V
167 723 208 0 1 3
0 12
0
0 0 54256 602
3 10V
-11 -15 10 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
6 74LS47
187 469 212 0 14 29
0 24 23 22 21 26 27 11 10 5
6 7 8 9 28
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
8 Hex Key~
166 307 165 0 11 12
0 20 19 18 17 0 0 0 0 0
1 49
0
0 0 4656 90
0
4 KPD2
-16 -27 12 -19
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7734 0 0
0
0
8 Hex Key~
166 306 201 0 11 12
0 16 15 14 13 0 0 0 0 0
1 49
0
0 0 4656 90
0
4 KPD1
-17 19 11 27
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9914 0 0
0
0
6 74LS83
105 382 186 0 14 29
0 20 19 18 17 16 15 14 13 2
24 23 22 21 3
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
9 Resistor~
219 695 206 0 4 5
0 4 12 0 1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
23
14 1 3 0 0 4240 0 8 1 0 0 3
414 231
414 289
415 289
1 9 2 0 0 4224 0 2 8 0 0 2
351 231
350 231
9 1 4 0 0 12416 0 3 9 0 0 5
555 69
555 65
669 65
669 206
677 206
9 5 5 0 0 8320 0 5 3 0 0 3
507 194
558 194
558 141
4 10 6 0 0 4224 0 3 5 0 0 3
552 141
552 203
507 203
3 11 7 0 0 4224 0 3 5 0 0 3
546 141
546 212
507 212
2 12 8 0 0 4224 0 3 5 0 0 3
540 141
540 221
507 221
1 13 9 0 0 4224 0 3 5 0 0 3
534 141
534 230
507 230
6 8 10 0 0 8320 0 3 5 0 0 3
564 141
564 185
507 185
7 7 11 0 0 8320 0 3 5 0 0 3
570 141
570 176
507 176
1 2 12 0 0 4224 0 4 9 0 0 2
712 206
713 206
4 8 13 0 0 4224 0 7 8 0 0 4
331 209
342 209
342 213
350 213
3 7 14 0 0 4224 0 7 8 0 0 4
331 203
342 203
342 204
350 204
2 6 15 0 0 4224 0 7 8 0 0 4
331 197
342 197
342 195
350 195
1 5 16 0 0 4224 0 7 8 0 0 4
331 191
342 191
342 186
350 186
4 4 17 0 0 4224 0 6 8 0 0 4
332 173
342 173
342 177
350 177
3 3 18 0 0 4224 0 6 8 0 0 4
332 167
342 167
342 168
350 168
2 2 19 0 0 4224 0 6 8 0 0 4
332 161
342 161
342 159
350 159
1 1 20 0 0 4224 0 6 8 0 0 4
332 155
342 155
342 150
350 150
4 13 21 0 0 4224 0 5 8 0 0 4
437 203
422 203
422 204
414 204
3 12 22 0 0 4224 0 5 8 0 0 4
437 194
422 194
422 195
414 195
2 11 23 0 0 4224 0 5 8 0 0 4
437 185
422 185
422 186
414 186
1 10 24 0 0 4224 0 5 8 0 0 4
437 176
422 176
422 177
414 177
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
