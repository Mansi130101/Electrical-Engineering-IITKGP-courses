CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 120 9
205 99 1280 689
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
205 99 1280 689
143654930 0
0
6 Title:
5 Name:
0
0
0
20
9 CA 7-Seg~
184 155 147 0 18 19
10 30 29 28 27 26 25 24 45 32
2 2 0 0 2 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8953 0 0
0
0
2 +V
167 155 50 0 1 3
0 31
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
6 74LS47
187 143 242 0 14 29
0 23 22 21 19 46 47 24 25 26
27 28 29 30 48
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3618 0 0
0
0
6 74LS93
109 177 324 0 8 17
0 2 2 20 19 23 22 21 19
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
7 Ground~
168 184 380 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Pulser~
4 64 378 0 10 12
0 49 50 20 51 0 0 5 5 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7734 0 0
0
0
7 Pulser~
4 384 385 0 10 12
0 52 53 5 54 0 0 5 5 3
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 504 387 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
6 74LS93
109 497 331 0 8 17
0 2 2 5 55 9 8 7 6
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U3
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
6 74LS47
187 463 249 0 14 29
0 9 8 7 6 56 57 10 11 12
13 14 15 16 58
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
2 +V
167 475 57 0 1 3
0 17
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
9 CA 7-Seg~
184 475 154 0 18 19
10 16 15 14 13 12 11 10 59 18
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8903 0 0
0
0
9 CA 7-Seg~
184 794 157 0 18 19
10 42 41 40 39 38 37 36 60 44
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3834 0 0
0
0
2 +V
167 794 60 0 1 3
0 43
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
6 74LS47
187 782 252 0 14 29
0 4 35 3 33 61 62 36 37 38
39 40 41 42 63
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U6
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
6 74LS93
109 816 334 0 8 17
0 4 3 34 33 4 35 3 33
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U5
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
7 Pulser~
4 703 388 0 10 12
0 64 65 34 66 0 0 5 5 3
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3874 0 0
0
0
9 Resistor~
219 155 85 0 4 5
0 32 31 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 475 92 0 4 5
0 18 17 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 794 95 0 4 5
0 44 43 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
50
2 3 3 0 0 12416 0 16 15 0 0 5
814 364
814 373
865 373
865 289
805 289
1 5 4 0 0 8320 0 16 16 0 0 4
823 364
862 364
862 300
823 300
3 3 5 0 0 4240 0 7 9 0 0 4
408 376
485 376
485 367
486 367
2 0 2 0 0 4112 0 9 0 0 5 3
495 361
495 376
504 376
1 1 2 0 0 4240 0 8 9 0 0 2
504 381
504 361
8 4 6 0 0 4240 0 9 10 0 0 2
477 297
477 286
7 3 7 0 0 4240 0 9 10 0 0 2
486 297
486 286
6 2 8 0 0 4240 0 9 10 0 0 2
495 297
495 286
5 1 9 0 0 4240 0 9 10 0 0 2
504 297
504 286
7 7 10 0 0 4240 0 10 12 0 0 4
504 216
504 196
490 196
490 190
8 6 11 0 0 4240 0 10 12 0 0 4
495 216
495 199
484 199
484 190
9 5 12 0 0 12432 0 10 12 0 0 4
486 216
486 204
478 204
478 190
10 4 13 0 0 12432 0 10 12 0 0 4
477 216
477 209
472 209
472 190
11 3 14 0 0 4240 0 10 12 0 0 4
468 216
468 198
466 198
466 190
12 2 15 0 0 4240 0 10 12 0 0 4
459 216
459 197
460 197
460 190
13 1 16 0 0 4240 0 10 12 0 0 4
450 216
450 198
454 198
454 190
1 2 17 0 0 4240 0 11 19 0 0 2
475 66
475 74
1 9 18 0 0 4240 0 19 12 0 0 2
475 110
475 118
4 0 19 0 0 12432 0 4 0 0 23 5
157 360
157 364
142 364
142 285
157 285
3 3 20 0 0 4240 0 6 4 0 0 4
88 369
165 369
165 360
166 360
2 0 2 0 0 16 0 4 0 0 22 3
175 354
175 369
184 369
1 1 2 0 0 16 0 5 4 0 0 2
184 374
184 354
8 4 19 0 0 16 0 4 3 0 0 2
157 290
157 279
7 3 21 0 0 4240 0 4 3 0 0 2
166 290
166 279
6 2 22 0 0 4240 0 4 3 0 0 2
175 290
175 279
5 1 23 0 0 4240 0 4 3 0 0 2
184 290
184 279
7 7 24 0 0 4240 0 3 1 0 0 4
184 209
184 189
170 189
170 183
8 6 25 0 0 4240 0 3 1 0 0 4
175 209
175 192
164 192
164 183
9 5 26 0 0 12432 0 3 1 0 0 4
166 209
166 197
158 197
158 183
10 4 27 0 0 12432 0 3 1 0 0 4
157 209
157 202
152 202
152 183
11 3 28 0 0 4240 0 3 1 0 0 4
148 209
148 191
146 191
146 183
12 2 29 0 0 4240 0 3 1 0 0 4
139 209
139 190
140 190
140 183
13 1 30 0 0 4240 0 3 1 0 0 4
130 209
130 191
134 191
134 183
1 2 31 0 0 4240 0 2 18 0 0 2
155 59
155 67
1 9 32 0 0 4240 0 18 1 0 0 2
155 103
155 111
4 0 33 0 0 12416 0 16 0 0 38 5
796 370
796 374
781 374
781 295
796 295
3 3 34 0 0 4224 0 17 16 0 0 4
727 379
804 379
804 370
805 370
8 4 33 0 0 0 0 16 15 0 0 2
796 300
796 289
7 3 3 0 0 0 0 16 15 0 0 2
805 300
805 289
6 2 35 0 0 4224 0 16 15 0 0 2
814 300
814 289
5 1 4 0 0 0 0 16 15 0 0 2
823 300
823 289
7 7 36 0 0 4224 0 15 13 0 0 4
823 219
823 199
809 199
809 193
8 6 37 0 0 4224 0 15 13 0 0 4
814 219
814 202
803 202
803 193
9 5 38 0 0 12416 0 15 13 0 0 4
805 219
805 207
797 207
797 193
10 4 39 0 0 12416 0 15 13 0 0 4
796 219
796 212
791 212
791 193
11 3 40 0 0 4224 0 15 13 0 0 4
787 219
787 201
785 201
785 193
12 2 41 0 0 4224 0 15 13 0 0 4
778 219
778 200
779 200
779 193
13 1 42 0 0 4224 0 15 13 0 0 4
769 219
769 201
773 201
773 193
1 2 43 0 0 4224 0 14 20 0 0 2
794 69
794 77
1 9 44 0 0 4224 0 20 13 0 0 2
794 113
794 121
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
0 1 2
0
0 0 100 100 0 0
77 66 1007 216
0 0 0 0
1007 66
77 66
1007 66
1007 216
0 0
5e-006 0 5e-006 0 5e-006 5e-006
12385 0
0 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
