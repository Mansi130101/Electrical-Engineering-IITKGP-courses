CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
340 0 20 80 9
402 83 1215 692
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
402 83 1215 692
177209362 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 213 526 0 1 11
0 3
0
0 0 21360 0
2 0V
-29 0 -15 8
2 V4
-31 -14 -17 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 172 472 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
14 12 28 20
2 V3
17 3 31 11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
7 Ground~
168 315 326 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 347 424 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 233 581 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
6 74LS47
187 768 501 0 14 29
0 14 15 16 17 48 49 10 9 8
7 6 5 4 50
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
3 U10
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
9 CA 7-Seg~
184 1093 317 0 17 19
10 4 5 6 7 8 9 10 51 42
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP8
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9914 0 0
0
0
9 Inverter~
13 1072 255 0 2 22
0 22 42
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 4 0
1 U
3747 0 0
0
0
9 CA 7-Seg~
184 1005 318 0 17 19
10 4 5 6 7 8 9 10 52 43
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP7
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
9 Inverter~
13 984 264 0 2 22
0 23 43
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
7931 0 0
0
0
9 Inverter~
13 888 273 0 2 22
0 24 44
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
9325 0 0
0
0
9 CA 7-Seg~
184 909 333 0 17 19
10 4 5 6 7 8 9 10 53 44
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8903 0 0
0
0
9 Inverter~
13 799 282 0 2 22
0 25 45
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 3 0
1 U
3834 0 0
0
0
9 CA 7-Seg~
184 820 335 0 17 19
10 4 5 6 7 8 9 10 54 45
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3363 0 0
0
0
9 Inverter~
13 707 291 0 2 22
0 26 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 3 0
1 U
7668 0 0
0
0
9 CA 7-Seg~
184 727 343 0 18 19
10 4 5 6 7 8 9 10 55 46
2 2 2 0 0 0 0 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4718 0 0
0
0
9 Inverter~
13 613 300 0 2 22
0 27 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 3 0
1 U
3874 0 0
0
0
9 CA 7-Seg~
184 634 344 0 17 19
10 4 5 6 7 8 9 10 56 11
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
6671 0 0
0
0
9 Inverter~
13 521 309 0 2 22
0 28 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 3 0
1 U
3789 0 0
0
0
9 CA 7-Seg~
184 542 362 0 17 19
10 4 5 6 7 8 9 10 57 12
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4871 0 0
0
0
9 CA 7-Seg~
184 450 359 0 17 19
10 4 5 6 7 8 9 10 58 13
2 2 2 0 0 0 0 2
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3750 0 0
0
0
7 74LS138
19 352 282 0 14 29
0 20 19 18 21 2 2 22 23 24
25 26 27 28 29
0
0 0 13296 0
7 74LS138
-26 58 23 66
2 U8
-6 49 8 57
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
9 Inverter~
13 429 318 0 2 22
0 29 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
538 0 0
0
0
10 Ascii Key~
169 580 543 0 11 12
0 33 32 31 30 59 60 61 36 0
0 57
0
0 0 4656 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
6843 0 0
0
0
7 74LS374
66 490 528 0 37 37
0 62 63 64 65 30 31 32 33 66
67 68 69 14 15 16 17 34 35 0
0 0 0 0 0 0 0 0 0 0
2 2 2 2 1 0 0 1
0
0 0 13040 512
7 74LS374
-24 -60 25 -52
2 U7
-13 -61 1 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 512 1 0 0 0
1 U
3136 0 0
0
0
7 74LS193
137 271 527 0 14 29
0 39 21 21 3 2 2 2 2 70
71 72 20 19 18
0
0 0 13040 0
7 74LS193
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5950 0 0
0
0
6 1K RAM
79 380 518 0 20 41
0 2 2 2 2 2 2 73 20 19
18 74 75 76 77 14 15 16 17 2
40
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U5
-7 57 7 65
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 0 0 0 0
1 U
5670 0 0
0
0
9 Inverter~
13 184 181 0 2 22
0 36 35
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
6828 0 0
0
0
7 Buffer~
58 142 181 0 2 22
0 35 37
0
0 0 624 512
4 4050
-14 -19 14 -11
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 2 0
1 U
6735 0 0
0
0
7 Buffer~
58 99 180 0 2 22
0 37 38
0
0 0 624 512
4 4050
-14 -19 14 -11
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 2 0
1 U
8365 0 0
0
0
5 4073~
219 81 249 0 4 22
0 38 37 35 34
0
0 0 624 0
6 74LS11
-14 -24 28 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
4132 0 0
0
0
7 Ground~
168 168 390 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4551 0 0
0
0
7 74LS157
122 131 432 0 14 29
0 47 41 34 78 79 21 34 80 81
2 39 82 40 83
0
0 0 13040 180
7 74LS157
-24 -60 25 -52
2 U1
-13 -61 1 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
3635 0 0
0
0
7 Pulser~
4 41 349 0 10 12
0 84 85 41 86 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3973 0 0
0
0
2 +V
167 51 431 0 1 3
0 21
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3851 0 0
0
0
123
19 1 2 0 0 8336 0 27 4 0 0 4
418 482
418 446
347 446
347 432
1 4 3 0 0 8320 0 1 26 0 0 3
225 526
225 527
239 527
8 7 2 0 0 0 0 26 26 0 0 2
239 563
239 554
1 8 2 0 0 0 0 5 26 0 0 3
233 575
233 563
239 563
1 0 2 0 0 0 0 3 0 0 75 2
315 320
314 318
1 10 2 0 0 0 0 32 33 0 0 2
161 391
163 391
1 0 2 0 0 0 0 4 0 0 111 3
347 432
348 434
348 482
13 0 4 0 0 4096 0 6 0 0 66 4
755 468
755 411
756 411
756 406
12 0 5 0 0 4096 0 6 0 0 59 4
764 468
764 416
765 416
765 411
11 0 6 0 0 4096 0 6 0 0 52 4
773 468
773 423
774 423
774 417
10 0 7 0 0 4096 0 6 0 0 45 2
782 468
782 425
9 0 8 0 0 4096 0 6 0 0 38 2
791 468
791 431
8 0 9 0 0 4096 0 6 0 0 31 4
800 468
800 444
801 444
801 439
7 0 10 0 0 4096 0 6 0 0 24 4
809 468
809 450
810 450
810 445
7 0 10 0 0 4096 0 9 0 0 24 4
1020 354
1020 440
1021 440
1021 445
7 0 10 0 0 0 0 12 0 0 24 2
924 369
924 445
7 0 10 0 0 0 0 14 0 0 24 4
835 371
835 440
836 440
836 445
7 0 10 0 0 0 0 16 0 0 24 2
742 379
742 445
7 0 10 0 0 0 0 18 0 0 24 2
649 380
649 445
7 0 10 0 0 0 0 20 0 0 24 2
557 398
557 445
2 9 11 0 0 4224 0 17 18 0 0 2
634 300
634 308
2 9 12 0 0 4224 0 19 20 0 0 2
542 309
542 326
2 9 13 0 0 4224 0 23 21 0 0 2
450 318
450 323
7 7 10 0 0 8320 0 21 7 0 0 4
465 395
465 445
1108 445
1108 353
6 0 9 0 0 8192 0 9 0 0 31 3
1014 354
1015 354
1015 439
6 0 9 0 0 0 0 12 0 0 31 2
918 369
918 439
6 0 9 0 0 0 0 14 0 0 31 2
829 371
829 439
6 0 9 0 0 0 0 16 0 0 31 3
736 379
736 439
737 439
6 0 9 0 0 0 0 18 0 0 31 3
643 380
644 380
644 439
6 0 9 0 0 0 0 20 0 0 31 2
551 398
551 439
6 6 9 0 0 8320 0 21 7 0 0 4
459 395
459 439
1102 439
1102 353
5 0 8 0 0 4096 0 9 0 0 38 2
1008 354
1008 431
5 0 8 0 0 0 0 12 0 0 38 4
912 369
912 393
913 393
913 431
5 0 8 0 0 0 0 14 0 0 38 2
823 371
823 431
5 0 8 0 0 0 0 16 0 0 38 4
730 379
730 434
731 434
731 431
5 0 8 0 0 0 0 18 0 0 38 4
637 380
637 434
638 434
638 431
5 0 8 0 0 0 0 20 0 0 38 2
545 398
545 431
5 5 8 0 0 8320 0 21 7 0 0 4
453 395
453 431
1096 431
1096 353
4 0 7 0 0 4096 0 9 0 0 45 2
1002 354
1002 425
4 0 7 0 0 0 0 12 0 0 45 2
906 369
906 425
4 0 7 0 0 0 0 14 0 0 45 2
817 371
817 425
4 0 7 0 0 0 0 16 0 0 45 3
724 379
725 379
725 425
4 0 7 0 0 0 0 18 0 0 45 5
631 380
633 380
633 394
632 394
632 425
4 0 7 0 0 0 0 20 0 0 45 2
539 398
539 425
4 4 7 0 0 8320 0 21 7 0 0 4
447 395
447 425
1090 425
1090 353
3 0 6 0 0 4096 0 9 0 0 52 2
996 354
996 417
3 0 6 0 0 0 0 12 0 0 52 2
900 369
900 417
3 0 6 0 0 0 0 14 0 0 52 3
811 371
812 371
812 417
3 0 6 0 0 0 0 16 0 0 52 3
718 379
719 379
719 417
3 0 6 0 0 0 0 18 0 0 52 3
625 380
626 380
626 417
3 0 6 0 0 0 0 20 0 0 52 3
533 398
532 398
532 417
3 3 6 0 0 8320 0 21 7 0 0 4
441 395
441 417
1084 417
1084 353
2 0 5 0 0 4096 0 9 0 0 59 2
990 354
990 411
2 0 5 0 0 0 0 12 0 0 59 2
894 369
894 411
2 0 5 0 0 0 0 14 0 0 59 2
805 371
805 411
2 0 5 0 0 0 0 18 0 0 59 3
619 380
620 380
620 411
2 0 5 0 0 0 0 20 0 0 59 3
527 398
526 398
526 411
2 0 5 0 0 0 0 16 0 0 59 4
712 379
712 393
713 393
713 411
2 2 5 0 0 8320 0 21 7 0 0 4
435 395
435 411
1078 411
1078 353
1 0 4 0 0 0 0 9 0 0 66 2
984 354
984 406
1 0 4 0 0 0 0 12 0 0 66 4
888 369
888 392
887 392
887 406
1 0 4 0 0 0 0 14 0 0 66 2
799 371
799 406
1 0 4 0 0 0 0 20 0 0 66 4
521 398
521 399
510 399
510 406
1 0 4 0 0 0 0 18 0 0 66 4
613 380
613 395
612 395
612 406
1 0 4 0 0 0 0 16 0 0 66 2
706 379
706 406
1 1 4 0 0 8320 0 21 7 0 0 4
429 395
429 406
1072 406
1072 353
1 13 14 0 0 8320 0 6 25 0 0 7
809 538
809 627
526 627
526 628
428 628
428 537
452 537
2 14 15 0 0 8320 0 6 25 0 0 5
800 538
800 616
432 616
432 546
452 546
3 15 16 0 0 8320 0 6 25 0 0 5
791 538
791 605
438 605
438 555
452 555
4 16 17 0 0 8320 0 6 25 0 0 5
782 538
782 594
444 594
444 564
452 564
3 0 18 0 0 8320 0 22 0 0 100 6
320 273
294 273
294 452
315 452
315 563
340 563
2 0 19 0 0 8320 0 22 0 0 101 7
320 264
301 264
301 445
324 445
324 553
334 553
334 554
1 0 20 0 0 8320 0 22 0 0 102 7
320 255
310 255
310 439
332 439
332 544
330 544
330 543
4 0 21 0 0 8192 0 22 0 0 104 4
320 300
241 300
241 441
216 441
5 6 2 0 0 0 0 22 22 0 0 2
314 309
314 318
7 1 22 0 0 4224 0 22 8 0 0 2
390 255
1057 255
8 1 23 0 0 4224 0 22 10 0 0 2
390 264
969 264
9 1 24 0 0 4224 0 22 11 0 0 2
390 273
873 273
10 1 25 0 0 4224 0 22 13 0 0 2
390 282
784 282
11 1 26 0 0 4224 0 22 15 0 0 2
390 291
692 291
12 1 27 0 0 4224 0 22 17 0 0 2
390 300
598 300
13 1 28 0 0 4224 0 22 19 0 0 2
390 309
506 309
14 1 29 0 0 4224 0 22 23 0 0 2
390 318
414 318
5 4 30 0 0 4224 0 25 24 0 0 4
516 537
548 537
548 546
556 546
6 3 31 0 0 12416 0 25 24 0 0 4
516 546
535 546
535 552
556 552
7 2 32 0 0 12416 0 25 24 0 0 4
516 555
529 555
529 558
556 558
8 1 33 0 0 4224 0 25 24 0 0 2
516 564
556 564
17 4 34 0 0 16512 0 25 31 0 0 7
522 492
522 470
491 470
491 224
177 224
177 249
102 249
18 1 35 0 0 20608 0 25 29 0 0 8
452 492
434 492
434 438
404 438
404 200
165 200
165 181
157 181
1 8 36 0 0 4224 0 28 24 0 0 6
205 181
582 181
582 472
548 472
548 522
556 522
1 3 35 0 0 0 0 29 31 0 0 6
157 181
161 181
161 119
25 119
25 258
57 258
1 2 37 0 0 16512 0 30 31 0 0 6
114 180
118 180
118 142
35 142
35 249
57 249
2 1 38 0 0 8320 0 30 31 0 0 4
84 180
49 180
49 240
57 240
2 1 35 0 0 0 0 28 29 0 0 2
169 181
157 181
2 1 37 0 0 0 0 29 30 0 0 4
127 181
122 181
122 180
114 180
18 16 17 0 0 0 0 27 25 0 0 4
412 563
444 563
444 564
452 564
17 15 16 0 0 0 0 27 25 0 0 4
412 554
444 554
444 555
452 555
16 14 15 0 0 0 0 27 25 0 0 4
412 545
444 545
444 546
452 546
15 13 14 0 0 0 0 27 25 0 0 4
412 536
444 536
444 537
452 537
14 10 18 0 0 0 0 26 27 0 0 6
303 563
340 563
340 562
340 562
340 563
348 563
13 9 19 0 0 0 0 26 27 0 0 2
303 554
348 554
12 8 20 0 0 0 0 26 27 0 0 6
303 545
330 545
330 543
340 543
340 545
348 545
2 3 21 0 0 0 0 26 26 0 0 4
239 509
218 509
218 518
233 518
3 1 21 0 0 12288 0 26 35 0 0 5
233 518
216 518
216 441
51 441
51 440
6 7 2 0 0 0 0 26 26 0 0 2
239 545
239 554
5 6 2 0 0 0 0 26 26 0 0 2
239 536
239 545
6 5 2 0 0 0 0 27 27 0 0 2
348 527
348 518
5 4 2 0 0 0 0 27 27 0 0 2
348 518
348 509
4 3 2 0 0 0 0 27 27 0 0 2
348 509
348 500
2 3 2 0 0 0 0 27 27 0 0 2
348 491
348 500
1 2 2 0 0 0 0 27 27 0 0 2
348 482
348 491
11 1 39 0 0 12416 0 33 26 0 0 4
93 454
85 454
85 500
239 500
13 20 40 0 0 12416 0 33 27 0 0 6
93 418
66 418
66 599
423 599
423 491
418 491
7 4 34 0 0 0 0 33 31 0 0 4
157 418
178 418
178 249
102 249
3 4 34 0 0 0 0 33 31 0 0 4
157 454
188 454
188 249
102 249
6 1 21 0 0 12416 0 33 35 0 0 6
157 427
199 427
199 375
30 375
30 440
51 440
3 2 41 0 0 4224 0 34 33 0 0 4
65 340
204 340
204 463
157 463
9 2 42 0 0 4224 0 7 8 0 0 2
1093 281
1093 255
9 2 43 0 0 4224 0 9 10 0 0 2
1005 282
1005 264
9 2 44 0 0 4224 0 12 11 0 0 2
909 297
909 273
9 2 45 0 0 4224 0 14 13 0 0 2
820 299
820 282
9 2 46 0 0 12416 0 16 15 0 0 4
727 307
727 306
728 306
728 291
1 1 47 0 0 4224 0 2 33 0 0 2
160 472
157 472
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
644 81 806 104
656 91 810 106
22 19ee10039 mansi uniyal
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
