CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 80 9
4 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
4 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
37
7 Ground~
168 625 826 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
6 74LS83
105 534 773 0 14 29
0 2 2 2 2 5 6 7 8 4
12 11 10 9 65
0
0 0 13040 602
7 74LS83A
-24 -60 25 -52
3 U15
56 -3 77 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4441 0 0
0
0
9 Inverter~
13 927 659 0 2 22
0 16 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
3618 0 0
0
0
8 2-In OR~
219 902 900 0 3 22
0 14 13 17
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U12A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6153 0 0
0
0
9 2-In AND~
219 921 952 0 3 22
0 15 17 35
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U13C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
5394 0 0
0
0
9 Inverter~
13 364 610 0 2 22
0 4 29
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 737 845 0 3 22
0 4 20 31
0
0 0 624 180
6 74LS86
-21 -24 21 -16
4 U14C
-5 -25 23 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 7 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 742 945 0 3 22
0 18 4 33
0
0 0 624 512
6 74LS86
-21 -24 21 -16
4 U14A
-5 -25 23 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 736 795 0 3 22
0 21 4 30
0
0 0 624 512
6 74LS86
-21 -24 21 -16
4 U14D
-5 -25 23 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 7 0
1 U
3549 0 0
0
0
9 2-In XOR~
219 741 894 0 3 22
0 19 4 32
0
0 0 624 512
6 74LS86
-21 -24 21 -16
4 U14B
-5 -25 23 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
7931 0 0
0
0
9 2-In AND~
219 838 632 0 3 22
0 34 16 4
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9325 0 0
0
0
9 Inverter~
13 870 643 0 2 22
0 13 34
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U11B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
8903 0 0
0
0
5 7405~
219 334 754 0 2 22
0 35 36
0
0 0 624 90
6 74LS05
-21 -24 21 -16
3 U9A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
3834 0 0
0
0
7 Ground~
168 636 873 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Ground~
168 973 848 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
7 74LS157
122 541 859 0 14 29
0 35 41 33 40 32 39 31 38 30
2 8 7 6 5
0
0 0 13040 90
7 74LS157
-24 -60 25 -52
3 U10
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
7 Ground~
168 1208 776 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
2 +V
167 1265 819 0 1 3
0 37
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6671 0 0
0
0
6 74LS83
105 1044 870 0 14 29
0 2 37 37 2 21 20 19 18 2
38 39 40 41 14
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
10 Ascii Key~
169 1116 40 0 11 12
0 64 63 62 61 66 67 68 60 0
0 54
0
0 0 4656 512
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
4871 0 0
0
0
7 74LS273
150 1140 164 0 18 37
0 3 55 69 70 71 72 61 62 63
64 73 74 75 76 43 44 45 46
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
7 74LS273
150 1140 282 0 18 37
0 3 55 77 78 79 80 43 44 45
46 81 82 83 84 56 16 57 58
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U3
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
6 74LS83
105 1035 688 0 14 29
0 51 52 53 54 47 48 49 50 16
21 20 19 18 13
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
6 74LS47
187 504 707 0 14 29
0 12 11 10 9 85 86 22 23 24
25 26 27 28 87
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6843 0 0
0
0
2 +V
167 1305 122 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3136 0 0
0
0
7 Buffer~
58 1137 96 0 2 22
0 60 55
0
0 0 624 270
4 4050
-14 -19 14 -11
3 U1A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
5950 0 0
0
0
2 +V
167 513 196 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5670 0 0
0
0
9 CA 7-Seg~
184 511 520 0 18 19
10 28 27 26 25 24 23 22 88 59
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6828 0 0
0
0
7 74LS273
150 1140 415 0 18 37
0 3 55 89 90 91 92 56 16 57
58 93 94 95 96 47 48 49 50
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U6
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
6735 0 0
0
0
9 2-In XOR~
219 1280 506 0 3 22
0 46 16 54
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
8365 0 0
0
0
9 2-In XOR~
219 1352 504 0 3 22
0 45 16 53
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
4132 0 0
0
0
9 2-In XOR~
219 1415 505 0 3 22
0 44 16 52
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
4551 0 0
0
0
9 2-In XOR~
219 1472 505 0 3 22
0 43 16 51
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3635 0 0
0
0
9 CA 7-Seg~
184 353 526 0 18 19
10 97 36 36 98 99 100 29 101 42
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3973 0 0
0
0
2 +V
167 355 202 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3851 0 0
0
0
9 Resistor~
219 512 281 0 4 5
0 59 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 356 272 0 4 5
0 42 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
101
9 0 4 0 0 8192 0 2 0 0 34 4
491 807
491 765
652 765
652 632
5 14 5 0 0 12432 0 2 16 0 0 5
536 807
541 807
541 816
572 816
572 826
13 6 6 0 0 4224 0 16 2 0 0 5
554 826
540 826
540 818
527 818
527 807
12 7 7 0 0 16512 0 16 2 0 0 5
536 826
528 826
528 820
518 820
518 807
11 8 8 0 0 12416 0 16 2 0 0 4
518 826
518 822
509 822
509 807
1 1 2 0 0 4096 0 2 1 0 0 3
572 807
625 807
625 820
2 1 2 0 0 0 0 2 2 0 0 2
563 807
572 807
3 2 2 0 0 0 0 2 2 0 0 2
554 807
563 807
4 3 2 0 0 0 0 2 2 0 0 2
545 807
554 807
13 4 9 0 0 4224 0 2 24 0 0 2
518 743
518 744
12 3 10 0 0 4224 0 2 24 0 0 2
527 743
527 744
11 2 11 0 0 4224 0 2 24 0 0 2
536 743
536 744
10 1 12 0 0 4224 0 2 24 0 0 2
545 743
545 744
2 0 13 0 0 4224 0 4 0 0 19 2
896 884
896 722
14 1 14 0 0 8320 0 19 4 0 0 3
1001 904
1001 884
914 884
2 1 15 0 0 4224 0 3 5 0 0 3
930 677
930 930
928 930
0 1 16 0 0 8192 0 0 3 41 0 3
931 623
930 623
930 641
3 2 17 0 0 4224 0 4 5 0 0 2
905 930
910 930
14 1 13 0 0 128 0 23 12 0 0 3
992 722
891 722
891 643
0 1 18 0 0 4224 0 0 8 59 0 4
1019 832
867 832
867 936
764 936
0 1 19 0 0 4224 0 0 10 58 0 4
1028 819
851 819
851 885
763 885
0 2 20 0 0 4224 0 0 7 57 0 4
1037 799
834 799
834 836
759 836
1 0 21 0 0 4224 0 9 0 0 56 2
758 786
1046 786
2 0 4 0 0 0 0 9 0 0 40 2
758 804
811 804
1 0 4 0 0 0 0 7 0 0 40 2
759 854
811 854
2 0 4 0 0 0 0 10 0 0 40 2
763 903
811 903
7 7 22 0 0 4224 0 28 24 0 0 4
526 556
526 624
545 624
545 674
6 8 23 0 0 4224 0 28 24 0 0 4
520 556
520 642
536 642
536 674
5 9 24 0 0 4224 0 28 24 0 0 4
514 556
514 650
527 650
527 674
4 10 25 0 0 4224 0 28 24 0 0 4
508 556
508 664
518 664
518 674
3 11 26 0 0 8320 0 28 24 0 0 5
502 556
503 556
503 671
509 671
509 674
2 12 27 0 0 8320 0 28 24 0 0 3
496 556
500 556
500 674
1 13 28 0 0 12416 0 28 24 0 0 4
490 556
490 571
491 571
491 674
3 1 4 0 0 4224 0 11 6 0 0 3
811 632
367 632
367 628
2 7 29 0 0 4224 0 6 34 0 0 3
367 592
367 562
368 562
3 9 30 0 0 8320 0 9 16 0 0 5
709 795
652 795
652 923
572 923
572 890
3 7 31 0 0 12416 0 7 16 0 0 5
710 845
681 845
681 939
554 939
554 890
3 5 32 0 0 12416 0 10 16 0 0 5
714 894
698 894
698 947
536 947
536 890
3 3 33 0 0 8320 0 16 8 0 0 4
518 890
518 960
715 960
715 945
3 2 4 0 0 128 0 11 8 0 0 3
811 632
811 954
764 954
2 0 16 0 0 4096 0 11 0 0 64 2
856 623
992 623
2 1 34 0 0 4224 0 12 11 0 0 3
855 643
855 641
856 641
10 1 2 0 0 0 0 16 14 0 0 4
581 896
581 908
629 908
629 874
1 0 35 0 0 8192 0 13 0 0 45 3
337 772
337 906
501 906
3 1 35 0 0 8320 0 5 16 0 0 6
919 975
919 971
501 971
501 906
500 906
500 890
3 0 36 0 0 4224 0 34 0 0 47 3
344 562
344 672
337 672
2 2 36 0 0 128 0 34 13 0 0 4
338 562
338 672
337 672
337 736
2 0 37 0 0 4096 0 19 0 0 49 3
1073 840
1073 836
1074 836
3 1 37 0 0 8320 0 19 18 0 0 4
1064 840
1064 836
1265 836
1265 828
1 1 2 0 0 8192 0 19 17 0 0 4
1082 840
1082 762
1208 762
1208 770
9 1 2 0 0 0 0 19 15 0 0 3
1001 840
1001 842
973 842
10 8 38 0 0 8320 0 19 16 0 0 4
1055 904
1055 1016
563 1016
563 890
11 6 39 0 0 8320 0 19 16 0 0 4
1046 904
1046 1005
545 1005
545 890
12 4 40 0 0 8320 0 19 16 0 0 4
1037 904
1037 996
527 996
527 890
2 13 41 0 0 8320 0 16 19 0 0 4
509 890
509 985
1028 985
1028 904
10 5 21 0 0 128 0 23 19 0 0 2
1046 722
1046 840
11 6 20 0 0 128 0 23 19 0 0 2
1037 722
1037 840
12 7 19 0 0 128 0 23 19 0 0 2
1028 722
1028 840
13 8 18 0 0 128 0 23 19 0 0 2
1019 722
1019 840
4 1 2 0 0 8320 0 19 17 0 0 4
1055 840
1055 759
1208 759
1208 770
9 0 42 0 0 4096 0 34 0 0 62 3
353 490
353 488
355 488
1 9 42 0 0 8320 0 37 0 0 61 4
356 290
355 290
355 490
353 490
2 1 3 0 0 4096 0 37 35 0 0 3
356 254
356 211
355 211
9 0 16 0 0 4224 0 23 0 0 82 3
992 658
992 332
1113 332
0 1 43 0 0 4224 0 0 33 94 0 3
1121 242
1484 242
1484 486
0 1 44 0 0 4224 0 0 32 95 0 3
1112 232
1427 232
1427 486
0 1 45 0 0 8320 0 0 31 96 0 3
1103 222
1364 222
1364 485
0 1 46 0 0 8320 0 0 30 97 0 3
1094 213
1292 213
1292 487
15 5 47 0 0 12416 0 29 23 0 0 4
1121 452
1121 495
1037 495
1037 658
16 6 48 0 0 12416 0 29 23 0 0 4
1112 452
1112 485
1028 485
1028 658
17 7 49 0 0 12416 0 29 23 0 0 4
1103 452
1103 475
1019 475
1019 658
18 8 50 0 0 12416 0 29 23 0 0 4
1094 452
1094 463
1010 463
1010 658
3 1 51 0 0 8320 0 33 23 0 0 4
1475 535
1475 568
1073 568
1073 658
3 2 52 0 0 8320 0 32 23 0 0 4
1418 535
1418 558
1064 558
1064 658
3 3 53 0 0 8320 0 31 23 0 0 4
1355 534
1355 547
1055 547
1055 658
3 4 54 0 0 8320 0 30 23 0 0 4
1283 536
1283 538
1046 538
1046 658
0 2 55 0 0 4224 0 0 29 87 0 4
1207 200
1207 368
1166 368
1166 388
0 1 3 0 0 4224 0 0 29 92 0 3
1220 249
1220 382
1175 382
0 2 16 0 0 0 0 0 33 80 0 3
1408 332
1466 332
1466 486
0 2 16 0 0 0 0 0 32 81 0 3
1341 332
1409 332
1409 486
0 2 16 0 0 0 0 0 31 82 0 3
1276 332
1346 332
1346 485
0 2 16 0 0 0 0 0 30 84 0 5
1113 332
1276 332
1276 332
1274 332
1274 487
15 7 56 0 0 4224 0 22 29 0 0 2
1121 319
1121 388
16 8 16 0 0 0 0 22 29 0 0 5
1112 319
1113 319
1113 332
1112 332
1112 388
17 9 57 0 0 4224 0 22 29 0 0 2
1103 319
1103 388
18 10 58 0 0 4224 0 22 29 0 0 2
1094 319
1094 388
0 2 55 0 0 0 0 0 22 88 0 6
1159 128
1159 116
1234 116
1234 200
1166 200
1166 255
2 2 55 0 0 0 0 26 21 0 0 4
1137 111
1137 128
1166 128
1166 137
1 9 59 0 0 4224 0 36 28 0 0 4
512 299
512 478
511 478
511 484
2 1 3 0 0 0 0 36 27 0 0 4
512 263
514 263
514 205
513 205
1 8 60 0 0 4224 0 26 20 0 0 2
1137 81
1137 64
1 1 3 0 0 0 0 22 25 0 0 3
1175 249
1305 249
1305 131
1 1 3 0 0 0 0 21 25 0 0 2
1175 131
1305 131
15 7 43 0 0 0 0 21 22 0 0 2
1121 201
1121 255
16 8 44 0 0 0 0 21 22 0 0 2
1112 201
1112 255
17 9 45 0 0 0 0 21 22 0 0 2
1103 201
1103 255
18 10 46 0 0 0 0 21 22 0 0 2
1094 201
1094 255
4 7 61 0 0 4224 0 20 21 0 0 4
1113 64
1113 130
1121 130
1121 137
3 8 62 0 0 4224 0 20 21 0 0 3
1107 64
1107 137
1112 137
2 9 63 0 0 8320 0 20 21 0 0 3
1101 64
1103 64
1103 137
1 10 64 0 0 8320 0 20 21 0 0 3
1095 64
1094 64
1094 137
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
1529 149 1615 191
1541 159 1619 189
23 MODI OMKAR 
19EE30018
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
0 0.05 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
