CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 70 1 80 9
638 79 1240 679
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
638 79 1240 679
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 545 107 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
8 2-In OR~
219 394 249 0 3 22
0 20 28 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 185696511
65 0 0 0 4 1 1 0
1 U
4441 0 0
0
0
9 8-In NOR~
219 384 330 0 9 19
0 27 26 25 24 23 22 21 28 20
0
0 0 624 90
4 4078
-7 -24 21 -16
2 U7
25 -1 39 7
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
7 Ground~
168 682 414 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 706 415 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Pulser~
4 637 158 0 10 12
0 50 51 30 52 0 0 5 5 6
7
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7734 0 0
0
0
2 +V
167 654 638 0 1 3
0 34
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
2 +V
167 899 618 0 1 3
0 35
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3747 0 0
0
0
9 CA 7-Seg~
184 822 684 0 18 19
10 42 41 40 39 38 37 36 53 32
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
9 CA 7-Seg~
184 618 684 0 18 19
10 49 48 47 46 45 44 43 54 33
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7931 0 0
0
0
6 74LS47
187 720 573 0 14 29
0 23 22 21 28 55 56 36 37 38
39 40 41 42 57
0
0 0 13040 270
7 74LS247
-24 -60 25 -52
2 U6
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
6 74LS47
187 529 578 0 14 29
0 27 26 25 24 58 59 43 44 45
46 47 48 49 60
0
0 0 13040 270
7 74LS247
-24 -60 25 -52
2 U5
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
6 74LS83
105 749 439 0 14 29
0 18 17 16 15 14 13 12 11 2
23 22 21 28 31
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
6 74LS83
105 559 438 0 14 29
0 3 4 5 6 7 8 9 10 31
27 26 25 24 61
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U3
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
7 74LS273
150 741 200 0 18 37
0 29 30 7 8 9 10 14 13 12
11 3 4 5 6 18 17 16 15
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
7 74LS273
150 543 201 0 18 37
0 29 30 27 26 25 24 23 22 21
19 7 8 9 10 14 13 12 11
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
9 Resistor~
219 636 647 0 4 5
0 33 34 0 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 880 627 0 4 5
0 32 35 0 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6671 0 0
0
0
76
1 11 3 0 0 8320 0 14 15 0 0 5
597 408
597 285
872 285
872 182
773 182
2 12 4 0 0 8320 0 14 15 0 0 5
588 408
588 291
868 291
868 191
773 191
3 13 5 0 0 8320 0 14 15 0 0 5
579 408
579 297
862 297
862 200
773 200
4 14 6 0 0 8320 0 14 15 0 0 5
570 408
570 307
855 307
855 209
773 209
5 0 7 0 0 4224 0 14 0 0 43 4
561 408
561 276
605 276
605 183
6 0 8 0 0 4224 0 14 0 0 44 4
552 408
552 272
600 272
600 192
7 0 9 0 0 4224 0 14 0 0 45 4
543 408
543 265
594 265
594 201
8 0 10 0 0 4224 0 14 0 0 46 4
534 408
534 260
586 260
586 210
8 0 11 0 0 12416 0 13 0 0 50 4
724 409
724 341
669 341
669 246
7 0 12 0 0 12416 0 13 0 0 49 4
733 409
733 337
679 337
679 237
6 0 13 0 0 12416 0 13 0 0 48 4
742 409
742 332
687 332
687 228
5 0 14 0 0 12416 0 13 0 0 47 4
751 409
751 327
694 327
694 219
4 18 15 0 0 4224 0 13 15 0 0 5
760 409
760 259
776 259
776 245
773 245
3 17 16 0 0 12416 0 13 15 0 0 7
769 409
769 346
787 346
787 259
788 259
788 236
773 236
2 16 17 0 0 12416 0 13 15 0 0 5
778 409
778 354
798 354
798 227
773 227
1 15 18 0 0 8320 0 13 15 0 0 4
787 409
827 409
827 218
773 218
3 10 19 0 0 8320 0 2 16 0 0 3
427 249
427 246
511 246
9 1 20 0 0 8320 0 3 2 0 0 4
390 297
355 297
355 240
381 240
7 0 21 0 0 8192 0 3 0 0 30 3
413 353
413 389
494 389
6 0 22 0 0 8192 0 3 0 0 28 3
404 353
404 399
485 399
5 0 23 0 0 8192 0 3 0 0 27 3
395 353
395 409
478 409
4 0 24 0 0 8192 0 3 0 0 31 3
386 353
386 435
470 435
3 0 25 0 0 8192 0 3 0 0 32 3
377 353
377 441
461 441
2 0 26 0 0 8192 0 3 0 0 33 3
368 353
368 450
451 450
1 0 27 0 0 8192 0 3 0 0 34 3
359 353
359 459
440 459
2 0 28 0 0 12288 0 2 0 0 29 7
381 258
370 258
370 289
434 289
434 354
426 354
426 352
0 7 23 0 0 8320 0 0 16 72 0 4
761 514
478 514
478 219
511 219
0 8 22 0 0 8320 0 0 16 71 0 4
752 521
485 521
485 228
511 228
4 8 28 0 0 12432 0 11 3 0 0 6
734 540
693 540
693 352
426 352
426 353
422 353
9 0 21 0 0 8320 0 16 0 0 70 4
511 237
494 237
494 529
743 529
0 6 24 0 0 8320 0 0 16 73 0 4
543 507
470 507
470 210
511 210
0 5 25 0 0 8320 0 0 16 74 0 4
552 501
461 501
461 201
511 201
0 4 26 0 0 8320 0 0 16 75 0 4
561 492
451 492
451 192
511 192
0 3 27 0 0 8320 0 0 16 76 0 4
570 484
440 484
440 183
511 183
1 1 29 0 0 8320 0 15 1 0 0 4
703 164
703 108
557 108
557 107
1 1 29 0 0 0 0 16 1 0 0 6
505 165
501 165
501 127
565 127
565 107
557 107
1 1 2 0 0 8320 0 5 4 0 0 4
706 409
706 400
682 400
682 408
1 9 2 0 0 0 0 5 13 0 0 2
706 409
706 409
2 3 30 0 0 12416 0 16 6 0 0 6
511 174
472 174
472 116
675 116
675 149
661 149
0 1 29 0 0 128 0 0 15 35 0 4
703 164
704 164
704 164
703 164
3 2 30 0 0 128 0 6 15 0 0 4
661 149
686 149
686 173
709 173
9 14 31 0 0 8320 0 14 13 0 0 6
516 408
516 449
664 449
664 481
706 481
706 473
11 3 7 0 0 0 0 16 15 0 0 4
575 183
695 183
695 182
709 182
12 4 8 0 0 0 0 16 15 0 0 4
575 192
695 192
695 191
709 191
13 5 9 0 0 0 0 16 15 0 0 4
575 201
695 201
695 200
709 200
14 6 10 0 0 0 0 16 15 0 0 4
575 210
695 210
695 209
709 209
15 7 14 0 0 0 0 16 15 0 0 4
575 219
695 219
695 218
709 218
16 8 13 0 0 0 0 16 15 0 0 4
575 228
695 228
695 227
709 227
17 9 12 0 0 0 0 16 15 0 0 4
575 237
695 237
695 236
709 236
18 10 11 0 0 0 0 16 15 0 0 4
575 246
695 246
695 245
709 245
9 1 32 0 0 8320 0 9 18 0 0 3
822 648
822 627
862 627
1 9 33 0 0 4224 0 17 10 0 0 2
618 647
618 648
2 1 34 0 0 0 0 17 7 0 0 2
654 647
654 647
2 1 35 0 0 4224 0 18 8 0 0 2
898 627
899 627
7 7 36 0 0 4224 0 11 9 0 0 4
761 610
761 728
837 728
837 720
8 6 37 0 0 4224 0 11 9 0 0 4
752 610
752 728
831 728
831 720
9 5 38 0 0 4224 0 11 9 0 0 4
743 610
743 728
825 728
825 720
10 4 39 0 0 4224 0 11 9 0 0 4
734 610
734 728
819 728
819 720
11 3 40 0 0 4224 0 11 9 0 0 4
725 610
725 728
813 728
813 720
12 2 41 0 0 4224 0 11 9 0 0 4
716 610
716 728
807 728
807 720
13 1 42 0 0 4224 0 11 9 0 0 4
707 610
707 728
801 728
801 720
7 7 43 0 0 4224 0 12 10 0 0 4
570 615
570 728
633 728
633 720
8 6 44 0 0 4224 0 12 10 0 0 4
561 615
561 728
627 728
627 720
9 5 45 0 0 4224 0 12 10 0 0 4
552 615
552 728
621 728
621 720
10 4 46 0 0 4224 0 12 10 0 0 4
543 615
543 728
615 728
615 720
11 3 47 0 0 4224 0 12 10 0 0 4
534 615
534 728
609 728
609 720
12 2 48 0 0 4224 0 12 10 0 0 4
525 615
525 728
603 728
603 720
13 1 49 0 0 4224 0 12 10 0 0 4
516 615
516 728
597 728
597 720
4 13 28 0 0 0 0 11 13 0 0 3
734 540
734 473
733 473
3 12 21 0 0 0 0 11 13 0 0 3
743 540
743 473
742 473
2 11 22 0 0 0 0 11 13 0 0 3
752 540
752 473
751 473
1 10 23 0 0 0 0 11 13 0 0 3
761 540
761 473
760 473
4 13 24 0 0 0 0 12 14 0 0 2
543 545
543 472
3 12 25 0 0 0 0 12 14 0 0 2
552 545
552 472
2 11 26 0 0 0 0 12 14 0 0 2
561 545
561 472
1 10 27 0 0 0 0 12 14 0 0 2
570 545
570 472
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
855 348 954 409
867 358 958 403
38 on the reset 
to start 
simulation
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
790 88 894 152
800 96 896 144
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
