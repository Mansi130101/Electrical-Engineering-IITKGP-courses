CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 80 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
143654930 0
0
6 Title:
5 Name:
0
0
0
37
2 +V
167 263 487 0 1 3
0 14
0
0 0 54256 0
2 5V
-19 -1 -5 7
2 V4
-5 -25 9 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 229 475 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 829 647 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
6 74LS83
105 804 570 0 14 29
0 4 5 6 7 2 2 2 2 25
24 23 22 3 3
0
0 0 13040 90
7 74LS83A
-24 -60 25 -52
3 U14
56 -3 77 5
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
7 Ground~
168 731 699 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
9 2-In XOR~
219 627 561 0 3 22
0 26 25 31
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U13D
-25 24 3 32
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 6 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 589 566 0 3 22
0 27 25 32
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U13C
-27 27 1 35
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 6 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 549 573 0 3 22
0 28 25 33
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U13B
-32 25 -4 33
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 6 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 503 578 0 3 22
0 29 25 34
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U13A
-26 29 2 37
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
3549 0 0
0
0
9 Inverter~
13 934 479 0 2 22
0 25 35
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 3 0
1 U
7931 0 0
0
0
9 Inverter~
13 903 462 0 2 22
0 8 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 3 0
1 U
9325 0 0
0
0
7 74LS157
122 691 655 0 14 29
0 8 9 34 10 33 11 32 12 31
2 7 6 5 4
0
0 0 13040 90
7 74LS157
-24 -60 25 -52
3 U12
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
8 2-In OR~
219 388 611 0 3 22
0 36 37 30
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U11A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1677489093
65 0 0 0 4 1 5 0
1 U
3834 0 0
0
0
9 2-In AND~
219 133 606 0 3 22
0 38 39 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U10B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
3363 0 0
0
0
9 Inverter~
13 119 567 0 2 22
0 36 39
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9B
-29 -5 -8 3
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
7668 0 0
0
0
9 2-In AND~
219 384 660 0 3 22
0 30 40 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U10A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1761375182
65 0 0 0 4 1 4 0
1 U
4718 0 0
0
0
9 Inverter~
13 381 476 0 2 22
0 38 40
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
3874 0 0
0
0
6 74LS83
105 269 534 0 14 29
0 26 27 28 29 2 14 14 2 2
12 11 10 9 37
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
2 +V
167 922 284 0 1 3
0 43
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V3
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
9 CA 7-Seg~
184 922 369 0 18 19
10 67 13 13 68 69 70 35 71 42
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
-42 -39 -7 -31
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4871 0 0
0
0
9 CA 7-Seg~
184 995 367 0 18 19
10 15 16 17 18 19 20 21 72 41
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-42 -39 -7 -31
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3750 0 0
0
0
2 +V
167 995 284 0 1 3
0 44
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8778 0 0
0
0
9 2-In XOR~
219 120 350 0 3 22
0 38 47 52
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7D
-23 29 -2 37
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
538 0 0
0
0
9 2-In XOR~
219 166 345 0 3 22
0 38 48 53
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7C
-29 25 -8 33
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6843 0 0
0
0
9 2-In XOR~
219 206 338 0 3 22
0 38 49 54
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7B
-24 27 -3 35
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3136 0 0
0
0
9 2-In XOR~
219 244 333 0 3 22
0 38 50 51
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7A
-22 24 -1 32
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1316181930
65 0 0 0 4 1 2 0
1 U
5950 0 0
0
0
7 74LS273
150 353 342 0 18 37
0 46 45 73 74 75 76 57 38 56
55 77 78 79 80 61 60 59 58
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
6 74LS83
105 296 417 0 14 29
0 61 60 59 58 51 54 53 52 38
26 27 28 29 36
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6828 0 0
0
0
14 Logic Display~
6 210 432 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
6 74LS47
187 1029 528 0 14 29
0 24 23 22 3 81 82 21 20 19
18 17 16 15 83
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8365 0 0
0
0
7 74LS273
150 353 266 0 18 37
0 46 45 84 85 86 87 50 49 48
47 88 89 90 91 57 38 56 55
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U6
53 13 67 21
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
4132 0 0
0
0
2 +V
167 440 108 0 1 3
0 46
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4551 0 0
0
0
10 Ascii Key~
169 330 48 0 11 12
0 66 65 64 63 92 93 94 62 0
0 56
0
0 0 4656 512
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3635 0 0
0
0
7 Buffer~
58 351 87 0 2 22
0 62 45
0
0 0 624 270
4 4050
-14 -19 14 -11
3 U3A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3973 0 0
0
0
7 74LS273
150 352 156 0 18 37
0 46 45 95 96 97 98 63 64 65
66 99 100 101 102 50 49 48 47
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3851 0 0
0
0
9 Resistor~
219 922 315 0 4 5
0 42 43 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 995 314 0 4 5
0 41 44 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
103
14 0 3 0 0 4096 0 4 0 0 23 2
847 540
847 534
14 1 4 0 0 8320 0 12 4 0 0 3
722 622
722 604
766 604
13 2 5 0 0 8320 0 12 4 0 0 4
704 622
704 609
775 609
775 604
12 3 6 0 0 8336 0 12 4 0 0 4
686 622
686 614
784 614
784 604
11 4 7 0 0 8320 0 12 4 0 0 4
668 622
668 617
793 617
793 604
0 1 8 0 0 12416 0 0 11 48 0 4
649 748
649 747
906 747
906 480
13 2 9 0 0 8320 0 18 12 0 0 4
253 568
253 740
659 740
659 686
12 4 10 0 0 8320 0 18 12 0 0 4
262 568
262 734
677 734
677 686
11 6 11 0 0 8320 0 18 12 0 0 4
271 568
271 728
695 728
695 686
10 8 12 0 0 8320 0 18 12 0 0 4
280 568
280 721
713 721
713 686
3 0 13 0 0 4096 0 20 0 0 12 3
913 405
913 413
907 413
2 2 13 0 0 4224 0 11 20 0 0 4
906 444
906 413
907 413
907 405
1 0 14 0 0 0 0 1 0 0 57 2
263 496
263 496
1 0 2 0 0 0 0 2 0 0 56 2
236 476
236 476
9 0 2 0 0 4096 0 18 0 0 56 2
226 504
236 504
13 1 15 0 0 4224 0 30 21 0 0 4
1048 495
1048 411
974 411
974 403
12 2 16 0 0 4224 0 30 21 0 0 4
1039 495
1039 411
980 411
980 403
11 3 17 0 0 4224 0 30 21 0 0 4
1030 495
1030 411
986 411
986 403
10 4 18 0 0 4224 0 30 21 0 0 4
1021 495
1021 411
992 411
992 403
9 5 19 0 0 4224 0 30 21 0 0 4
1012 495
1012 411
998 411
998 403
8 6 20 0 0 4224 0 30 21 0 0 4
1003 495
1003 411
1004 411
1004 403
7 7 21 0 0 4224 0 30 21 0 0 4
994 495
994 411
1010 411
1010 403
13 4 3 0 0 8320 0 4 30 0 0 6
820 540
820 534
956 534
956 598
1021 598
1021 565
12 3 22 0 0 8320 0 4 30 0 0 6
811 540
811 530
960 530
960 592
1012 592
1012 565
11 2 23 0 0 8320 0 4 30 0 0 6
802 540
802 525
966 525
966 585
1003 585
1003 565
10 1 24 0 0 8320 0 4 30 0 0 6
793 540
793 521
974 521
974 573
994 573
994 565
5 6 2 0 0 0 0 4 4 0 0 2
802 604
811 604
7 6 2 0 0 0 0 4 4 0 0 2
820 604
811 604
1 7 2 0 0 8192 0 3 4 0 0 4
829 641
830 641
830 604
820 604
1 8 2 0 0 4224 0 3 4 0 0 4
829 641
829 595
829 595
829 604
9 0 25 0 0 4096 0 4 0 0 47 2
847 604
847 755
0 1 26 0 0 4224 0 0 6 62 0 3
307 504
639 504
639 542
0 1 27 0 0 12416 0 0 7 61 0 5
298 495
370 495
370 509
601 509
601 547
0 1 28 0 0 12416 0 0 8 60 0 5
289 484
370 484
370 514
561 514
561 554
0 1 29 0 0 12416 0 0 9 59 0 5
280 474
370 474
370 520
515 520
515 559
1 3 30 0 0 4224 0 16 13 0 0 2
391 638
391 641
3 9 31 0 0 4224 0 6 12 0 0 4
630 591
630 692
722 692
722 686
3 7 32 0 0 8320 0 7 12 0 0 4
592 596
592 699
704 699
704 686
3 5 33 0 0 8320 0 8 12 0 0 4
552 603
552 705
686 705
686 686
3 3 34 0 0 8320 0 9 12 0 0 4
506 608
506 711
668 711
668 686
1 10 2 0 0 0 0 5 12 0 0 2
731 693
731 692
0 2 25 0 0 0 0 0 6 43 0 4
583 534
583 529
621 529
621 542
0 2 25 0 0 0 0 0 7 44 0 4
543 541
543 534
583 534
583 547
0 2 25 0 0 0 0 0 8 45 0 4
497 546
497 541
543 541
543 554
0 2 25 0 0 4096 0 0 9 47 0 5
131 629
337 629
337 546
497 546
497 559
2 7 35 0 0 4224 0 10 20 0 0 2
937 461
937 405
3 1 25 0 0 8320 0 14 10 0 0 4
131 629
131 755
937 755
937 497
3 1 8 0 0 0 0 16 12 0 0 5
382 683
382 748
649 748
649 686
650 686
0 1 36 0 0 8320 0 0 13 53 0 4
165 449
165 530
400 530
400 595
14 2 37 0 0 8320 0 18 13 0 0 4
226 568
226 580
382 580
382 595
0 1 38 0 0 8192 0 0 14 73 0 3
239 456
140 456
140 584
2 2 39 0 0 4224 0 14 15 0 0 2
122 584
122 585
1 1 36 0 0 0 0 29 15 0 0 4
210 450
210 449
122 449
122 549
2 2 40 0 0 12416 0 17 16 0 0 5
384 494
384 499
359 499
359 638
373 638
1 0 38 0 0 0 0 17 0 0 73 2
384 458
384 459
5 8 2 0 0 128 0 18 18 0 0 5
271 504
271 476
236 476
236 504
244 504
0 0 14 0 0 8320 0 0 0 0 58 3
253 497
253 496
263 496
6 7 14 0 0 0 0 18 18 0 0 5
262 504
263 504
263 496
253 496
253 504
4 13 29 0 0 0 0 18 28 0 0 2
280 504
280 451
3 12 28 0 0 0 0 18 28 0 0 2
289 504
289 451
2 11 27 0 0 0 0 18 28 0 0 2
298 504
298 451
1 10 26 0 0 0 0 18 28 0 0 2
307 504
307 451
1 9 41 0 0 4224 0 37 21 0 0 2
995 332
995 331
1 9 42 0 0 4224 0 36 20 0 0 4
922 333
922 332
922 332
922 333
1 2 43 0 0 4224 0 19 36 0 0 2
922 293
922 297
1 2 44 0 0 4224 0 22 37 0 0 2
995 293
995 296
2 0 45 0 0 8320 0 27 0 0 92 3
379 315
424 315
424 186
0 1 46 0 0 4096 0 0 27 93 0 4
440 227
440 301
388 301
388 309
2 0 47 0 0 8320 0 23 0 0 100 3
114 331
114 229
307 229
2 0 48 0 0 8320 0 24 0 0 101 3
160 326
160 221
316 221
2 0 49 0 0 8320 0 25 0 0 102 3
200 319
200 210
325 210
2 15 50 0 0 4224 0 26 35 0 0 4
238 314
238 201
333 201
333 193
9 0 38 0 0 16512 0 28 0 0 74 8
253 387
253 384
239 384
239 459
463 459
463 288
325 288
325 306
0 0 38 0 0 0 0 0 0 75 84 4
255 298
255 287
325 287
325 306
0 1 38 0 0 0 0 0 26 76 0 4
218 297
218 298
256 298
256 314
0 1 38 0 0 0 0 0 25 77 0 3
177 297
218 297
218 319
1 1 38 0 0 0 0 23 24 0 0 4
132 331
132 297
178 297
178 326
3 5 51 0 0 4224 0 26 28 0 0 3
247 363
298 363
298 387
3 8 52 0 0 4224 0 23 28 0 0 3
123 380
271 380
271 387
3 7 53 0 0 4224 0 24 28 0 0 3
169 375
280 375
280 387
3 6 54 0 0 8320 0 25 28 0 0 4
209 368
209 369
289 369
289 387
10 18 55 0 0 4224 0 27 31 0 0 2
307 315
307 303
9 17 56 0 0 4224 0 27 31 0 0 2
316 315
316 303
8 16 38 0 0 0 0 27 31 0 0 2
325 315
325 303
7 15 57 0 0 4224 0 27 31 0 0 2
334 315
334 303
18 4 58 0 0 12416 0 27 28 0 0 4
307 379
307 378
307 378
307 387
17 3 59 0 0 12416 0 27 28 0 0 4
316 379
316 378
316 378
316 387
16 2 60 0 0 12416 0 27 28 0 0 4
325 379
325 378
325 378
325 387
15 1 61 0 0 12416 0 27 28 0 0 4
334 379
334 378
334 378
334 387
1 14 36 0 0 0 0 29 28 0 0 3
210 450
253 450
253 451
1 8 62 0 0 0 0 34 33 0 0 2
351 72
351 72
2 0 45 0 0 0 0 31 0 0 95 8
379 239
379 193
424 193
424 104
378 104
378 111
378 111
378 103
1 1 46 0 0 4224 0 32 31 0 0 4
440 117
440 229
388 229
388 233
1 1 46 0 0 0 0 35 32 0 0 4
387 123
387 119
440 119
440 117
2 2 45 0 0 0 0 35 34 0 0 4
378 129
378 103
351 103
351 102
4 7 63 0 0 4224 0 33 35 0 0 4
327 72
327 115
333 115
333 129
3 8 64 0 0 4224 0 33 35 0 0 4
321 72
321 115
324 115
324 129
2 9 65 0 0 4224 0 33 35 0 0 2
315 72
315 129
1 10 66 0 0 4224 0 33 35 0 0 4
309 72
309 115
306 115
306 129
10 18 47 0 0 0 0 31 35 0 0 3
307 239
307 193
306 193
9 17 48 0 0 0 0 31 35 0 0 3
316 239
316 193
315 193
8 16 49 0 0 0 0 31 35 0 0 3
325 239
325 193
324 193
7 15 50 0 0 0 0 31 35 0 0 3
334 239
334 193
333 193
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 310
489 171 736 403
501 181 740 361
310 Decimal 2 digit display calculator

1. default tens digit blank (all 
low)
2. when negative only g high all 
low
3. if addition>9 and <15, +6 and 
display, tens digit displays 1
4. if addition>15 carry 1 +6 add 
and tens display 1
5. if subtraction negative (carry 
0) then display g(-ve sign).
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
