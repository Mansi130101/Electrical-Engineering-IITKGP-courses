CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
1 80 1281 689
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 80 1281 689
143654930 0
0
6 Title:
5 Name:
0
0
0
5
6 74LS47
187 212 250 0 14 29
0 2 12 13 14 15 16 3 4 5
6 7 8 9 17
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8953 0 0
0
0
7 Ground~
168 253 302 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
2 +V
167 224 58 0 1 3
0 10
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
9 CA 7-Seg~
184 224 155 0 18 19
10 9 8 7 6 5 4 3 18 11
0 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
6153 0 0
0
0
9 Resistor~
219 224 93 0 4 5
0 11 10 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
10
1 1 2 0 0 4224 0 2 1 0 0 2
253 296
253 287
7 7 3 0 0 4224 0 1 4 0 0 4
253 217
253 197
239 197
239 191
8 6 4 0 0 4224 0 1 4 0 0 4
244 217
244 200
233 200
233 191
9 5 5 0 0 12432 0 1 4 0 0 4
235 217
235 205
227 205
227 191
10 4 6 0 0 12416 0 1 4 0 0 4
226 217
226 210
221 210
221 191
11 3 7 0 0 4224 0 1 4 0 0 4
217 217
217 199
215 199
215 191
12 2 8 0 0 4224 0 1 4 0 0 4
208 217
208 198
209 198
209 191
13 1 9 0 0 4224 0 1 4 0 0 4
199 217
199 199
203 199
203 191
1 2 10 0 0 4224 0 3 5 0 0 2
224 67
224 75
1 9 11 0 0 4224 0 5 4 0 0 2
224 111
224 119
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
347 196 427 217
355 203 427 218
9 code 0111
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
