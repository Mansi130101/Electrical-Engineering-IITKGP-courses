CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 9
-9 79 775 688
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-9 79 775 688
143654930 0
0
6 Title:
5 Name:
0
0
0
16
9 2-In XOR~
219 120 350 0 3 22
0 8 4 11
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7D
-23 29 -2 37
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
8953 0 0
0
0
9 2-In XOR~
219 166 345 0 3 22
0 8 5 12
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7C
-29 25 -8 33
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
4441 0 0
0
0
9 2-In XOR~
219 206 338 0 3 22
0 8 6 13
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7B
-24 27 -3 35
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3618 0 0
0
0
9 2-In XOR~
219 244 333 0 3 22
0 8 7 10
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7A
-22 24 -1 32
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1316181930
65 0 0 0 4 1 2 0
1 U
6153 0 0
0
0
7 74LS273
150 353 342 0 18 37
0 3 2 39 40 41 42 20 8 19
18 43 44 45 46 24 23 22 21
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
6 74LS83
105 296 417 0 14 29
0 24 23 22 21 10 13 12 11 8
17 16 15 14 32
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7734 0 0
0
0
9 CA 7-Seg~
184 149 500 0 18 19
10 25 26 27 28 30 29 31 47 33
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-62 -24 -27 -16
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9914 0 0
0
0
2 +V
167 149 417 0 1 3
0 9
0
0 0 54256 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
14 Logic Display~
6 222 432 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
6 74LS47
187 267 497 0 14 29
0 17 16 15 14 48 49 31 29 30
28 27 26 25 50
0
0 0 13040 270
6 74LS47
-21 -60 21 -52
2 U1
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 74LS273
150 353 266 0 18 37
0 3 2 51 52 53 54 7 6 5
4 55 56 57 58 20 8 19 18
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U6
53 13 67 21
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
2 +V
167 440 108 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
10 Ascii Key~
169 330 48 0 11 12
0 38 37 36 35 59 60 61 34 0
0 57
0
0 0 4656 512
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3834 0 0
0
0
7 Buffer~
58 351 87 0 2 22
0 34 2
0
0 0 624 270
4 4050
-14 -19 14 -11
3 U3A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3363 0 0
0
0
7 74LS273
150 352 156 0 18 37
0 3 2 62 63 64 65 35 36 37
38 66 67 68 69 7 6 5 4
0
0 0 13040 270
7 74LS273
-24 -60 25 -52
2 U2
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
9 Resistor~
219 149 444 0 4 5
0 33 9 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
50
2 0 2 0 0 8336 0 5 0 0 39 3
379 315
424 315
424 186
0 1 3 0 0 4096 0 0 5 40 0 4
440 227
440 301
388 301
388 309
2 0 4 0 0 8320 0 1 0 0 47 3
114 331
114 229
307 229
2 0 5 0 0 8320 0 2 0 0 48 3
160 326
160 221
316 221
2 0 6 0 0 8320 0 3 0 0 49 3
200 319
200 210
325 210
2 15 7 0 0 4224 0 4 15 0 0 4
238 314
238 201
333 201
333 193
9 0 8 0 0 16512 0 6 0 0 8 8
253 387
253 384
239 384
239 455
463 455
463 288
325 288
325 306
0 0 8 0 0 0 0 0 0 9 23 4
255 298
255 256
325 256
325 306
0 1 8 0 0 0 0 0 4 11 0 4
218 297
218 298
256 298
256 314
1 2 9 0 0 0 0 8 16 0 0 2
149 426
149 426
0 1 8 0 0 0 0 0 3 12 0 3
177 297
218 297
218 319
1 1 8 0 0 0 0 1 2 0 0 4
132 331
132 297
178 297
178 326
3 5 10 0 0 4224 0 4 6 0 0 3
247 363
298 363
298 387
3 8 11 0 0 4224 0 1 6 0 0 3
123 380
271 380
271 387
3 7 12 0 0 4224 0 2 6 0 0 3
169 375
280 375
280 387
3 6 13 0 0 8320 0 3 6 0 0 4
209 368
209 369
289 369
289 387
4 13 14 0 0 4224 0 10 6 0 0 3
281 464
281 451
280 451
3 12 15 0 0 4224 0 10 6 0 0 3
290 464
290 451
289 451
2 11 16 0 0 4224 0 10 6 0 0 3
299 464
299 451
298 451
1 10 17 0 0 4224 0 10 6 0 0 3
308 464
308 451
307 451
10 18 18 0 0 4224 0 5 11 0 0 2
307 315
307 303
9 17 19 0 0 4224 0 5 11 0 0 2
316 315
316 303
8 16 8 0 0 128 0 5 11 0 0 2
325 315
325 303
7 15 20 0 0 4224 0 5 11 0 0 2
334 315
334 303
18 4 21 0 0 12416 0 5 6 0 0 4
307 379
307 378
307 378
307 387
17 3 22 0 0 12416 0 5 6 0 0 4
316 379
316 378
316 378
316 387
16 2 23 0 0 12416 0 5 6 0 0 4
325 379
325 378
325 378
325 387
15 1 24 0 0 12416 0 5 6 0 0 4
334 379
334 378
334 378
334 387
13 1 25 0 0 8320 0 10 7 0 0 4
254 534
254 620
128 620
128 536
2 12 26 0 0 8320 0 7 10 0 0 4
134 536
134 598
263 598
263 534
3 11 27 0 0 8320 0 7 10 0 0 4
140 536
140 589
272 589
272 534
4 10 28 0 0 8320 0 7 10 0 0 4
146 536
146 579
281 579
281 534
6 8 29 0 0 8320 0 7 10 0 0 4
158 536
158 557
299 557
299 534
5 9 30 0 0 8320 0 7 10 0 0 4
152 536
152 566
290 566
290 534
7 7 31 0 0 8320 0 7 10 0 0 4
164 536
164 545
308 545
308 534
1 14 32 0 0 4224 0 9 6 0 0 3
222 450
253 450
253 451
1 9 33 0 0 12416 0 16 7 0 0 4
149 462
149 442
149 442
149 464
1 8 34 0 0 0 0 14 13 0 0 2
351 72
351 72
2 0 2 0 0 128 0 11 0 0 42 8
379 239
379 193
424 193
424 104
378 104
378 111
378 111
378 103
1 1 3 0 0 4224 0 12 11 0 0 4
440 117
440 229
388 229
388 233
1 1 3 0 0 0 0 15 12 0 0 4
387 123
387 119
440 119
440 117
2 2 2 0 0 0 0 15 14 0 0 4
378 129
378 103
351 103
351 102
4 7 35 0 0 4224 0 13 15 0 0 4
327 72
327 115
333 115
333 129
3 8 36 0 0 4224 0 13 15 0 0 4
321 72
321 115
324 115
324 129
2 9 37 0 0 4224 0 13 15 0 0 2
315 72
315 129
1 10 38 0 0 4224 0 13 15 0 0 4
309 72
309 115
306 115
306 129
10 18 4 0 0 0 0 11 15 0 0 3
307 239
307 193
306 193
9 17 5 0 0 0 0 11 15 0 0 3
316 239
316 193
315 193
8 16 6 0 0 0 0 11 15 0 0 3
325 239
325 193
324 193
7 15 7 0 0 0 0 11 15 0 0 3
334 239
334 193
333 193
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 169
520 171 738 289
532 181 742 271
169 single digit calculator using 
3 74273 to memorize the 
operand (+/-) and using the 
XOR for the case of 
subtraction to generate 1s 
compliment of the number.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
