CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
430 110 5 80 9
638 79 1240 679
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
638 79 1240 679
143654930 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 662 408 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
2 +V
167 704 156 0 1 3
0 2
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
7 Pulser~
4 637 158 0 10 12
0 50 51 3 52 0 0 5 5 5
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3618 0 0
0
0
2 +V
167 504 156 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
7 Pulser~
4 462 183 0 10 12
0 53 54 4 55 0 0 5 5 5
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5394 0 0
0
0
2 +V
167 654 638 0 1 3
0 34
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
2 +V
167 899 618 0 1 3
0 35
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
9 CA 7-Seg~
184 822 684 0 18 19
10 42 41 40 39 38 37 36 56 32
2 0 2 2 2 0 0 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3747 0 0
0
0
9 CA 7-Seg~
184 618 684 0 18 19
10 49 48 47 46 45 44 43 57 33
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
6 74LS47
187 720 573 0 14 29
0 19 18 17 16 58 59 36 37 38
39 40 41 42 60
0
0 0 13040 270
7 74LS247
-24 -60 25 -52
2 U6
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
6 74LS47
187 529 578 0 14 29
0 23 22 21 20 61 62 43 44 45
46 47 48 49 63
0
0 0 13040 270
7 74LS247
-24 -60 25 -52
2 U5
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
6 74LS83
105 749 439 0 14 29
0 31 30 29 28 11 10 9 8 6
19 18 17 16 7
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
6 74LS83
105 559 438 0 14 29
0 27 26 25 24 15 14 13 12 7
23 22 21 20 64
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U3
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
7 74LS273
150 741 200 0 18 37
0 2 3 8 9 10 11 12 13 14
15 28 29 30 31 24 25 26 27
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
7 74LS273
150 543 201 0 18 37
0 5 4 16 17 18 19 20 21 22
23 8 9 10 11 12 13 14 15
0
0 0 13040 0
7 74LS273
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
9 Resistor~
219 636 647 0 4 5
0 33 34 0 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 880 627 0 4 5
0 32 35 0 1
0
0 0 880 0
3 330
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3874 0 0
0
0
64
1 1 2 0 0 4224 0 2 14 0 0 3
704 165
704 164
703 164
3 2 3 0 0 4224 0 3 14 0 0 4
661 149
686 149
686 173
709 173
3 2 4 0 0 4224 0 5 15 0 0 2
486 174
511 174
1 1 5 0 0 4224 0 4 15 0 0 2
504 165
505 165
1 9 6 0 0 8320 0 1 12 0 0 3
674 408
674 409
706 409
9 14 7 0 0 8320 0 13 12 0 0 6
516 408
516 449
691 449
691 481
706 481
706 473
11 3 8 0 0 4096 0 15 14 0 0 4
575 183
695 183
695 182
709 182
12 4 9 0 0 4096 0 15 14 0 0 4
575 192
695 192
695 191
709 191
13 5 10 0 0 4096 0 15 14 0 0 4
575 201
695 201
695 200
709 200
14 6 11 0 0 4096 0 15 14 0 0 4
575 210
695 210
695 209
709 209
15 7 12 0 0 4096 0 15 14 0 0 4
575 219
695 219
695 218
709 218
16 8 13 0 0 4096 0 15 14 0 0 4
575 228
695 228
695 227
709 227
17 9 14 0 0 4096 0 15 14 0 0 4
575 237
695 237
695 236
709 236
18 10 15 0 0 4096 0 15 14 0 0 4
575 246
695 246
695 245
709 245
3 0 16 0 0 8320 0 15 0 0 57 4
511 183
501 183
501 529
734 529
4 0 17 0 0 8320 0 15 0 0 58 4
511 192
501 192
501 523
743 523
5 0 18 0 0 8320 0 15 0 0 59 4
511 201
501 201
501 517
752 517
6 0 19 0 0 8320 0 15 0 0 60 4
511 210
501 210
501 511
761 511
7 0 20 0 0 8320 0 15 0 0 61 4
511 219
501 219
501 504
543 504
8 0 21 0 0 8320 0 15 0 0 62 4
511 228
501 228
501 498
552 498
9 0 22 0 0 8320 0 15 0 0 63 4
511 237
501 237
501 491
561 491
10 0 23 0 0 8320 0 15 0 0 64 4
511 246
501 246
501 483
570 483
4 15 24 0 0 8320 0 13 14 0 0 5
570 408
570 333
781 333
781 218
773 218
3 16 25 0 0 8320 0 13 14 0 0 5
579 408
579 324
781 324
781 227
773 227
2 17 26 0 0 8320 0 13 14 0 0 5
588 408
588 315
781 315
781 236
773 236
1 18 27 0 0 8320 0 13 14 0 0 5
597 408
597 309
781 309
781 245
773 245
4 11 28 0 0 12416 0 12 14 0 0 5
760 409
760 390
800 390
800 182
773 182
3 12 29 0 0 12416 0 12 14 0 0 5
769 409
769 397
811 397
811 191
773 191
2 13 30 0 0 12416 0 12 14 0 0 5
778 409
778 404
819 404
819 200
773 200
1 14 31 0 0 8320 0 12 14 0 0 4
787 409
828 409
828 209
773 209
8 3 8 0 0 12416 0 12 14 0 0 5
724 409
724 390
659 390
659 182
709 182
7 4 9 0 0 12416 0 12 14 0 0 5
733 409
733 382
670 382
670 191
709 191
6 5 10 0 0 12416 0 12 14 0 0 5
742 409
742 374
680 374
680 200
709 200
5 6 11 0 0 12416 0 12 14 0 0 5
751 409
751 369
688 369
688 209
709 209
8 15 12 0 0 4224 0 13 15 0 0 5
534 408
534 260
583 260
583 219
575 219
7 16 13 0 0 4224 0 13 15 0 0 5
543 408
543 260
583 260
583 228
575 228
6 17 14 0 0 4224 0 13 15 0 0 5
552 408
552 260
583 260
583 237
575 237
5 18 15 0 0 4224 0 13 15 0 0 5
561 408
561 260
583 260
583 246
575 246
9 1 32 0 0 8320 0 8 17 0 0 3
822 648
822 627
862 627
1 9 33 0 0 4224 0 16 9 0 0 2
618 647
618 648
2 1 34 0 0 0 0 16 6 0 0 2
654 647
654 647
2 1 35 0 0 4224 0 17 7 0 0 2
898 627
899 627
7 7 36 0 0 4224 0 10 8 0 0 4
761 610
761 728
837 728
837 720
8 6 37 0 0 4224 0 10 8 0 0 4
752 610
752 728
831 728
831 720
9 5 38 0 0 4224 0 10 8 0 0 4
743 610
743 728
825 728
825 720
10 4 39 0 0 4224 0 10 8 0 0 4
734 610
734 728
819 728
819 720
11 3 40 0 0 4224 0 10 8 0 0 4
725 610
725 728
813 728
813 720
12 2 41 0 0 4224 0 10 8 0 0 4
716 610
716 728
807 728
807 720
13 1 42 0 0 4224 0 10 8 0 0 4
707 610
707 728
801 728
801 720
7 7 43 0 0 4224 0 11 9 0 0 4
570 615
570 728
633 728
633 720
8 6 44 0 0 4224 0 11 9 0 0 4
561 615
561 728
627 728
627 720
9 5 45 0 0 4224 0 11 9 0 0 4
552 615
552 728
621 728
621 720
10 4 46 0 0 4224 0 11 9 0 0 4
543 615
543 728
615 728
615 720
11 3 47 0 0 4224 0 11 9 0 0 4
534 615
534 728
609 728
609 720
12 2 48 0 0 4224 0 11 9 0 0 4
525 615
525 728
603 728
603 720
13 1 49 0 0 4224 0 11 9 0 0 4
516 615
516 728
597 728
597 720
4 13 16 0 0 0 0 10 12 0 0 3
734 540
734 473
733 473
3 12 17 0 0 0 0 10 12 0 0 3
743 540
743 473
742 473
2 11 18 0 0 0 0 10 12 0 0 3
752 540
752 473
751 473
1 10 19 0 0 0 0 10 12 0 0 3
761 540
761 473
760 473
4 13 20 0 0 0 0 11 13 0 0 2
543 545
543 472
3 12 21 0 0 0 0 11 13 0 0 2
552 545
552 472
2 11 22 0 0 0 0 11 13 0 0 2
561 545
561 472
1 10 23 0 0 0 0 11 13 0 0 2
570 545
570 472
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
1026 187 1130 251
1036 195 1132 243
23 MANSI UNIYAL
19EE10039
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
