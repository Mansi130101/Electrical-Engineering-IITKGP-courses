CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 100 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
143654930 0
0
6 Title:
5 Name:
0
0
0
31
6 74LS93
109 870 335 0 8 17
0 4 5 3 6 4 7 5 6
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U9
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
8953 0 0
0
0
6 74LS47
187 836 253 0 14 29
0 4 7 5 6 62 63 8 9 10
11 12 13 14 64
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
3 U10
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4441 0 0
0
0
2 +V
167 848 61 0 1 3
0 15
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
9 CA 7-Seg~
184 848 158 0 18 19
10 14 13 12 11 10 9 8 65 16
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6153 0 0
0
0
8 2-In OR~
219 294 261 0 3 22
0 21 22 23
0
0 0 608 512
6 74LS32
-21 -24 21 -16
4 U12B
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
5394 0 0
0
0
8 2-In OR~
219 353 235 0 3 22
0 17 20 21
0
0 0 608 512
6 74LS32
-21 -24 21 -16
4 U12A
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 4 0
1 U
7734 0 0
0
0
8 2-In OR~
219 353 284 0 3 22
0 19 18 22
0
0 0 608 512
6 74LS32
-21 -24 21 -16
3 U2D
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -9401314
65 0 0 0 4 4 2 0
1 U
9914 0 0
0
0
8 2-In OR~
219 390 326 0 3 22
0 19 24 26
0
0 0 608 692
6 74LS32
-21 -24 21 -16
3 U2C
-37 -3 -16 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3747 0 0
0
0
9 2-In NOR~
219 237 352 0 3 22
0 23 25 24
0
0 0 608 602
6 74LS02
-21 -24 21 -16
4 U11A
-33 -20 -5 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -193950699
65 0 0 0 4 1 3 0
1 U
3549 0 0
0
0
8 2-In OR~
219 173 299 0 3 22
0 24 25 27
0
0 0 608 602
6 74LS32
-21 -24 21 -16
3 U2B
-35 -19 -14 -11
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -193950699
65 0 0 0 4 2 2 0
1 U
7931 0 0
0
0
8 2-In OR~
219 415 418 0 3 22
0 30 29 28
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 800149019
65 0 0 0 4 1 2 0
1 U
9325 0 0
0
0
9 2-In AND~
219 307 389 0 3 22
0 19 25 30
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
14 -13 35 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 1018187273
65 0 0 0 4 2 1 0
1 U
8903 0 0
0
0
9 2-In AND~
219 473 460 0 3 22
0 18 19 29
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U1A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 615599632
65 0 0 0 4 1 1 0
1 U
3834 0 0
0
0
7 Pulser~
4 805 394 0 10 12
0 66 67 3 68 0 0 5 5 6
7
0
0 0 4640 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3363 0 0
0
0
6 74LS93
109 649 340 0 8 17
0 40 50 4 51 52 40 50 51
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U6
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
6 74LS47
187 615 258 0 14 29
0 52 40 50 51 69 70 53 54 55
56 57 58 59 71
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
2 +V
167 627 66 0 1 3
0 60
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
9 CA 7-Seg~
184 627 163 0 18 19
10 59 58 57 56 55 54 53 72 61
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6671 0 0
0
0
6 74LS93
109 487 346 0 8 17
0 28 73 40 17 18 20 19 17
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U3
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
6 74LS47
187 453 244 0 14 29
0 18 20 26 17 74 75 41 42 43
44 45 46 47 76
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
2 +V
167 465 52 0 1 3
0 48
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3750 0 0
0
0
9 CA 7-Seg~
184 465 149 0 18 19
10 47 46 45 44 43 42 41 77 49
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8778 0 0
0
0
9 CA 7-Seg~
184 174 133 0 18 19
10 37 36 35 34 33 32 31 78 39
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
538 0 0
0
0
2 +V
167 174 41 0 1 3
0 38
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6843 0 0
0
0
6 74LS47
187 162 233 0 14 29
0 2 2 2 27 79 80 31 32 33
34 35 36 37 81
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3136 0 0
0
0
6 74LS93
109 187 382 0 8 17
0 30 82 29 25 83 84 85 25
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U8
27 3 41 11
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
5950 0 0
0
0
7 Ground~
168 242 276 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5670 0 0
0
0
9 Resistor~
219 848 96 0 4 5
0 16 15 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 627 101 0 4 5
0 61 60 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 465 87 0 4 5
0 49 48 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 174 76 0 4 5
0 39 38 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
84
3 3 3 0 0 4224 0 14 1 0 0 3
829 385
859 385
859 371
3 0 4 0 0 8320 0 15 0 0 4 4
638 376
638 422
895 422
895 373
2 0 5 0 0 12416 0 1 0 0 7 5
868 365
868 381
929 381
929 294
859 294
1 5 4 0 0 0 0 1 1 0 0 5
877 365
877 373
917 373
917 301
877 301
4 0 6 0 0 12416 0 1 0 0 6 5
850 371
850 375
835 375
835 301
850 301
8 4 6 0 0 0 0 1 2 0 0 2
850 301
850 290
7 3 5 0 0 0 0 1 2 0 0 2
859 301
859 290
6 2 7 0 0 4224 0 1 2 0 0 2
868 301
868 290
5 1 4 0 0 0 0 1 2 0 0 2
877 301
877 290
7 7 8 0 0 4224 0 2 4 0 0 4
877 220
877 200
863 200
863 194
8 6 9 0 0 4224 0 2 4 0 0 4
868 220
868 203
857 203
857 194
9 5 10 0 0 12416 0 2 4 0 0 4
859 220
859 208
851 208
851 194
10 4 11 0 0 12416 0 2 4 0 0 4
850 220
850 213
845 213
845 194
11 3 12 0 0 4224 0 2 4 0 0 4
841 220
841 202
839 202
839 194
12 2 13 0 0 4224 0 2 4 0 0 4
832 220
832 201
833 201
833 194
13 1 14 0 0 4224 0 2 4 0 0 4
823 220
823 202
827 202
827 194
1 2 15 0 0 4224 0 3 28 0 0 2
848 70
848 78
1 9 16 0 0 4224 0 28 4 0 0 2
848 114
848 122
4 1 17 0 0 8320 0 20 6 0 0 5
467 281
467 285
394 285
394 226
372 226
2 5 18 0 0 12288 0 7 19 0 0 5
372 293
376 293
376 299
494 299
494 312
1 7 19 0 0 12288 0 7 19 0 0 5
372 275
384 275
384 296
476 296
476 312
2 2 20 0 0 12416 0 6 20 0 0 5
372 244
389 244
389 292
485 292
485 281
2 7 19 0 0 8320 0 13 19 0 0 5
493 469
532 469
532 304
476 304
476 312
3 1 21 0 0 4224 0 6 5 0 0 3
326 235
326 252
313 252
3 2 22 0 0 4224 0 7 5 0 0 3
326 284
326 270
313 270
3 1 23 0 0 4224 0 5 9 0 0 4
267 261
267 385
252 385
252 371
2 3 24 0 0 4224 0 8 9 0 0 3
377 317
243 317
243 319
2 8 25 0 0 12288 0 9 26 0 0 5
234 371
222 371
222 345
167 345
167 348
1 3 24 0 0 0 0 10 9 0 0 4
185 315
185 317
243 317
243 319
1 7 19 0 0 0 0 8 19 0 0 7
377 335
371 335
371 347
432 347
432 302
476 302
476 312
3 3 26 0 0 8320 0 8 20 0 0 4
423 326
423 288
476 288
476 281
8 2 25 0 0 0 0 26 10 0 0 2
167 348
167 315
3 4 27 0 0 4224 0 10 25 0 0 2
176 269
176 270
7 1 19 0 0 0 0 19 12 0 0 6
476 312
476 306
440 306
440 368
283 368
283 380
2 8 25 0 0 8320 0 12 26 0 0 5
283 398
283 397
146 397
146 348
167 348
4 8 25 0 0 0 0 26 26 0 0 4
167 418
154 418
154 348
167 348
3 1 28 0 0 4224 0 11 19 0 0 3
448 418
494 418
494 376
2 0 29 0 0 8192 0 11 0 0 41 3
402 427
385 427
385 460
0 1 30 0 0 8192 0 0 11 40 0 3
334 410
334 409
402 409
3 1 30 0 0 12416 0 12 26 0 0 4
328 389
334 389
334 412
194 412
3 3 29 0 0 4224 0 13 26 0 0 3
448 460
176 460
176 418
5 1 18 0 0 8320 0 19 13 0 0 4
494 312
522 312
522 451
493 451
2 1 2 0 0 4096 0 25 25 0 0 2
194 270
203 270
2 3 2 0 0 0 0 25 25 0 0 2
194 270
185 270
1 1 2 0 0 4224 0 27 25 0 0 2
242 270
203 270
7 7 31 0 0 4224 0 25 23 0 0 4
203 200
203 180
189 180
189 169
8 6 32 0 0 4224 0 25 23 0 0 4
194 200
194 183
183 183
183 169
9 5 33 0 0 12416 0 25 23 0 0 4
185 200
185 188
177 188
177 169
10 4 34 0 0 12416 0 25 23 0 0 4
176 200
176 193
171 193
171 169
11 3 35 0 0 4224 0 25 23 0 0 4
167 200
167 182
165 182
165 169
12 2 36 0 0 4224 0 25 23 0 0 4
158 200
158 181
159 181
159 169
13 1 37 0 0 4224 0 25 23 0 0 4
149 200
149 182
153 182
153 169
1 2 38 0 0 4224 0 24 31 0 0 2
174 50
174 58
1 9 39 0 0 4224 0 31 23 0 0 4
174 94
174 98
174 98
174 97
0 3 40 0 0 12416 0 0 19 74 0 5
647 301
726 301
726 399
476 399
476 382
4 0 17 0 0 0 0 19 0 0 57 4
467 382
449 382
449 312
467 312
8 4 17 0 0 0 0 19 20 0 0 2
467 312
467 281
6 2 20 0 0 0 0 19 20 0 0 2
485 312
485 281
5 1 18 0 0 0 0 19 20 0 0 2
494 312
494 281
7 7 41 0 0 4224 0 20 22 0 0 4
494 211
494 191
480 191
480 185
8 6 42 0 0 4224 0 20 22 0 0 4
485 211
485 194
474 194
474 185
9 5 43 0 0 12416 0 20 22 0 0 4
476 211
476 199
468 199
468 185
10 4 44 0 0 12416 0 20 22 0 0 4
467 211
467 204
462 204
462 185
11 3 45 0 0 4224 0 20 22 0 0 4
458 211
458 193
456 193
456 185
12 2 46 0 0 4224 0 20 22 0 0 4
449 211
449 192
450 192
450 185
13 1 47 0 0 4224 0 20 22 0 0 4
440 211
440 193
444 193
444 185
1 2 48 0 0 4224 0 21 30 0 0 2
465 61
465 69
1 9 49 0 0 4224 0 30 22 0 0 2
465 105
465 113
2 3 50 0 0 12416 0 15 16 0 0 5
647 370
647 383
702 383
702 295
638 295
1 6 40 0 0 0 0 15 15 0 0 5
656 370
656 377
694 377
694 306
647 306
4 0 51 0 0 12416 0 15 0 0 72 5
629 376
629 380
614 380
614 306
629 306
8 4 51 0 0 0 0 15 16 0 0 2
629 306
629 295
7 3 50 0 0 0 0 15 16 0 0 2
638 306
638 295
6 2 40 0 0 0 0 15 16 0 0 2
647 306
647 295
5 1 52 0 0 4224 0 15 16 0 0 2
656 306
656 295
7 7 53 0 0 4224 0 16 18 0 0 4
656 225
656 205
642 205
642 199
8 6 54 0 0 4224 0 16 18 0 0 4
647 225
647 208
636 208
636 199
9 5 55 0 0 12416 0 16 18 0 0 4
638 225
638 213
630 213
630 199
10 4 56 0 0 12416 0 16 18 0 0 4
629 225
629 218
624 218
624 199
11 3 57 0 0 4224 0 16 18 0 0 4
620 225
620 207
618 207
618 199
12 2 58 0 0 4224 0 16 18 0 0 4
611 225
611 206
612 206
612 199
13 1 59 0 0 4224 0 16 18 0 0 4
602 225
602 207
606 207
606 199
1 2 60 0 0 4224 0 17 29 0 0 2
627 75
627 83
1 9 61 0 0 4224 0 29 18 0 0 2
627 119
627 127
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
1008 154 1120 198
1018 162 1122 194
25 MANSI UNIYAL 
19EE10039
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 196
959 199 1207 383
969 207 1209 351
196 Modifications on 24hr clock 
to make 12hr clock are:

1. minutes display remains 
the same
2. hours display resets at 12 
ie. modulo 12
3. converting 00 display on 
hours to 12 display
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
