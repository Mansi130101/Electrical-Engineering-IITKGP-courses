CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
420 50 30 120 9
0 71 1279 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1279 680
143654930 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 959 362 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 922 354 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
8 Hex Key~
166 762 361 0 11 12
0 5 4 3 2 0 0 0 0 0
9 57
0
0 0 4400 0
1 A
-3 -34 4 -26
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3618 0 0
0
0
8 Hex Key~
166 812 318 0 11 12
0 9 8 7 6 0 0 0 0 0
0 48
0
0 0 4400 0
1 S
-3 -34 4 -26
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6153 0 0
0
0
8 Hex Key~
166 703 391 0 11 12
0 13 10 11 12 0 0 0 0 0
6 54
0
0 0 4400 0
1 B
-3 -34 4 -26
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5394 0 0
0
0
14 Logic Display~
6 955 379 0 1 2
10 14
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L1
-2 15 12 23
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
12 Hex Display~
7 1009 400 0 18 19
10 15 16 17 18 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
2 0V
-8 -42 6 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9914 0 0
0
0
7 74LS181
132 879 399 0 22 45
0 6 7 8 9 2 3 4 5 12
11 10 13 20 19 14 21 22 23 18
17 16 15
0
0 0 13040 0
7 74LS181
-24 -69 25 -61
2 U8
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
19
4 5 2 0 0 8320 0 3 8 0 0 3
753 385
753 390
841 390
3 6 3 0 0 8320 0 3 8 0 0 3
759 385
759 399
841 399
2 7 4 0 0 8320 0 3 8 0 0 3
765 385
765 408
841 408
1 8 5 0 0 8320 0 3 8 0 0 3
771 385
771 417
841 417
4 1 6 0 0 8320 0 4 8 0 0 3
803 342
803 354
847 354
3 2 7 0 0 8320 0 4 8 0 0 3
809 342
809 363
847 363
2 3 8 0 0 8320 0 4 8 0 0 3
815 342
815 372
847 372
1 4 9 0 0 4224 0 4 8 0 0 3
821 342
821 381
847 381
2 11 10 0 0 8320 0 5 8 0 0 3
706 415
706 444
841 444
3 10 11 0 0 8320 0 5 8 0 0 3
700 415
700 435
841 435
4 9 12 0 0 8320 0 5 8 0 0 3
694 415
694 426
841 426
1 12 13 0 0 8320 0 5 8 0 0 3
712 415
712 453
841 453
1 15 14 0 0 8320 0 6 8 0 0 4
940 382
940 383
911 383
911 390
1 22 15 0 0 8320 0 7 8 0 0 3
1018 424
1018 453
917 453
2 21 16 0 0 8320 0 7 8 0 0 3
1012 424
1012 444
917 444
3 20 17 0 0 8320 0 7 8 0 0 3
1006 424
1006 435
917 435
4 19 18 0 0 8320 0 7 8 0 0 3
1000 424
1000 426
917 426
14 1 19 0 0 8320 0 8 1 0 0 3
911 363
911 362
947 362
1 13 20 0 0 4224 0 2 8 0 0 2
910 354
911 354
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
1026 187 1130 251
1036 195 1132 243
23 MANSI UNIYAL
19EE10039
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
1024 237 1165 336
1036 247 1169 322
51 74181 IC
A:9
B:Random generated 
other than 0,1
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
