CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 80 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
32
9 2-In NOR~
219 403 346 0 3 22
0 5 4 15
0
0 0 608 90
6 74LS02
-21 -24 21 -16
3 U7C
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -2034245009
65 0 0 0 4 3 1 0
1 U
8953 0 0
0
0
7 Ground~
168 420 297 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
4441 0 0
0
0
9 2-In AND~
219 551 488 0 3 22
0 10 6 9
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3618 0 0
0
0
9 Inverter~
13 538 534 0 2 22
0 7 10
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U10B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
6153 0 0
0
0
8 2-In OR~
219 577 451 0 3 22
0 9 5 8
0
0 0 608 692
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
5394 0 0
0
0
9 2-In AND~
219 719 447 0 3 22
0 11 7 12
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7734 0 0
0
0
9 Inverter~
13 706 508 0 2 22
0 6 11
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U10A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
9914 0 0
0
0
9 2-In AND~
219 495 396 0 3 22
0 6 7 4
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3747 0 0
0
0
9 2-In AND~
219 327 392 0 3 22
0 17 16 5
0
0 0 608 90
6 74LS08
-21 -24 21 -16
3 U8A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1950424477
65 0 0 0 4 1 2 0
1 U
3549 0 0
0
0
9 2-In NOR~
219 365 473 0 3 22
0 13 7 16
0
0 0 608 90
6 74LS02
-21 -24 21 -16
3 U7B
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
7931 0 0
0
0
9 2-In NOR~
219 271 472 0 3 22
0 14 6 17
0
0 0 608 90
6 74LS02
-21 -24 21 -16
3 U7A
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2051087763
65 0 0 0 4 1 1 0
1 U
9325 0 0
0
0
7 Ground~
168 996 388 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 1292 276 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
3834 0 0
0
0
2 +V
167 345 115 0 1 3
0 3
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V8
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
9 CA 7-Seg~
184 343 249 0 18 19
10 51 15 15 52 53 54 55 56 20
2 1 1 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7668 0 0
0
0
9 CA 7-Seg~
184 641 252 0 18 19
10 21 22 23 24 25 26 27 57 28
2 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4718 0 0
0
0
2 +V
167 643 118 0 1 3
0 3
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
6 74LS47
187 615 345 0 14 29
0 12 13 8 14 58 59 27 26 25
24 23 22 21 60
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
6 74LS93
109 648 679 0 8 17
0 7 13 18 14 7 13 6 14
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U6
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
9 CA 7-Seg~
184 918 252 0 18 19
10 31 32 33 34 35 36 37 61 38
2 0 0 2 2 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4871 0 0
0
0
2 +V
167 920 118 0 1 3
0 3
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3750 0 0
0
0
6 74LS47
187 892 345 0 14 29
0 2 18 29 30 62 63 37 36 35
34 33 32 31 64
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
6 74LS93
109 925 435 0 8 17
0 18 29 19 30 65 18 29 30
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U3
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
538 0 0
0
0
7 Pulser~
4 1071 520 0 10 12
0 66 67 41 68 0 0 5 5 4
7
0
0 0 4640 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6843 0 0
0
0
6 74LS93
109 1156 437 0 8 17
0 19 39 41 40 19 42 39 40
0
0 0 13024 602
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
6 74LS47
187 1124 349 0 14 29
0 19 42 39 40 69 70 49 48 47
46 45 44 43 71
0
0 0 13024 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5950 0 0
0
0
2 +V
167 1152 122 0 1 3
0 3
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5670 0 0
0
0
9 CA 7-Seg~
184 1150 256 0 18 19
10 43 44 45 46 47 48 49 72 50
0 0 0 0 2 2 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6828 0 0
0
0
9 Resistor~
219 344 169 0 4 5
0 20 3 0 1
0
0 0 864 90
3 330
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 642 172 0 4 5
0 28 3 0 1
0
0 0 864 90
3 330
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 919 172 0 4 5
0 38 3 0 1
0
0 0 864 90
3 330
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 1151 176 0 4 5
0 50 3 0 1
0
0 0 864 90
3 330
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
75
2 0 4 0 0 4096 0 1 0 0 19 2
418 365
419 365
1 0 5 0 0 4096 0 1 0 0 10 4
400 365
400 367
401 367
401 368
1 0 6 0 0 4096 0 8 0 0 25 2
485 417
485 601
2 0 7 0 0 4096 0 8 0 0 23 2
503 417
503 570
3 3 8 0 0 4224 0 18 5 0 0 3
638 382
638 451
610 451
1 3 9 0 0 4224 0 5 3 0 0 3
564 460
550 460
550 464
2 0 6 0 0 0 0 3 0 0 25 2
559 509
559 601
1 0 7 0 0 0 0 4 0 0 23 2
541 552
541 570
1 2 10 0 0 4224 0 3 4 0 0 2
541 509
541 516
0 2 5 0 0 8320 0 0 5 20 0 3
401 368
401 442
564 442
2 0 7 0 0 0 0 6 0 0 23 3
727 468
727 610
655 610
1 0 6 0 0 0 0 7 0 0 25 3
709 526
709 601
637 601
1 2 11 0 0 4224 0 6 7 0 0 2
709 468
709 490
1 3 12 0 0 8320 0 18 6 0 0 3
656 382
656 423
718 423
2 0 13 0 0 8192 0 18 0 0 24 3
647 382
646 382
646 585
4 0 14 0 0 8192 0 18 0 0 30 3
629 382
628 382
628 625
3 0 15 0 0 4096 0 15 0 0 18 2
334 285
334 316
2 3 15 0 0 8320 0 15 1 0 0 4
328 285
328 316
409 316
409 313
0 3 4 0 0 8320 0 0 8 0 0 4
419 362
419 367
494 367
494 372
3 0 5 0 0 0 0 9 0 0 0 3
326 368
401 368
401 362
3 2 16 0 0 8320 0 10 9 0 0 4
371 440
371 424
335 424
335 413
3 1 17 0 0 8320 0 11 9 0 0 4
277 439
277 424
317 424
317 413
2 5 7 0 0 8320 0 10 19 0 0 4
380 492
380 570
655 570
655 645
1 0 13 0 0 8320 0 10 0 0 29 4
362 492
362 582
646 582
646 622
2 7 6 0 0 8320 0 11 19 0 0 4
286 491
286 601
637 601
637 645
1 0 14 0 0 8320 0 11 0 0 30 3
268 491
268 622
584 622
1 1 2 0 0 4224 0 22 12 0 0 2
933 382
996 382
5 1 7 0 0 0 0 19 19 0 0 6
655 645
655 635
704 635
704 726
655 726
655 709
6 2 13 0 0 0 0 19 19 0 0 6
646 645
646 622
715 622
715 740
646 740
646 709
4 8 14 0 0 0 0 19 19 0 0 6
628 715
628 741
584 741
584 622
628 622
628 645
0 3 18 0 0 8320 0 0 19 49 0 5
924 387
978 387
978 787
637 787
637 715
0 1 18 0 0 0 0 0 23 49 0 6
924 399
924 395
951 395
951 495
932 495
932 465
1 3 19 0 0 12416 0 26 23 0 0 5
1165 386
1219 386
1219 587
914 587
914 471
1 2 3 0 0 4224 0 14 29 0 0 4
345 124
345 143
344 143
344 151
1 9 20 0 0 4224 0 29 15 0 0 4
344 187
344 205
343 205
343 213
1 13 21 0 0 8320 0 16 18 0 0 3
620 288
602 288
602 312
2 12 22 0 0 12416 0 16 18 0 0 4
626 288
626 293
611 293
611 312
3 11 23 0 0 12416 0 16 18 0 0 4
632 288
632 297
620 297
620 312
4 10 24 0 0 12416 0 16 18 0 0 4
638 288
638 299
629 299
629 312
5 9 25 0 0 8320 0 16 18 0 0 6
644 288
645 288
645 300
640 300
640 312
638 312
6 8 26 0 0 4224 0 16 18 0 0 3
650 288
650 312
647 312
7 7 27 0 0 4224 0 16 18 0 0 2
656 288
656 312
1 2 3 0 0 0 0 17 30 0 0 4
643 127
643 146
642 146
642 154
1 9 28 0 0 4224 0 30 16 0 0 4
642 190
642 208
641 208
641 216
0 2 29 0 0 8320 0 0 23 48 0 5
915 391
965 391
965 507
923 507
923 465
8 4 30 0 0 8320 0 23 23 0 0 5
905 401
873 401
873 473
905 473
905 471
8 4 30 0 0 0 0 23 22 0 0 3
905 401
906 401
906 382
7 3 29 0 0 0 0 23 22 0 0 3
914 401
915 401
915 382
6 2 18 0 0 0 0 23 22 0 0 3
923 401
924 401
924 382
1 13 31 0 0 8320 0 20 22 0 0 3
897 288
879 288
879 312
2 12 32 0 0 12416 0 20 22 0 0 4
903 288
903 293
888 293
888 312
3 11 33 0 0 12416 0 20 22 0 0 4
909 288
909 297
897 297
897 312
4 10 34 0 0 12416 0 20 22 0 0 4
915 288
915 299
906 299
906 312
5 9 35 0 0 8320 0 20 22 0 0 6
921 288
922 288
922 300
917 300
917 312
915 312
6 8 36 0 0 4224 0 20 22 0 0 3
927 288
927 312
924 312
7 7 37 0 0 4224 0 20 22 0 0 2
933 288
933 312
1 2 3 0 0 0 0 21 31 0 0 4
920 127
920 146
919 146
919 154
1 9 38 0 0 4224 0 31 20 0 0 4
919 190
919 208
918 208
918 216
0 1 19 0 0 0 0 0 25 66 0 7
1165 403
1183 403
1183 490
1164 490
1164 468
1163 468
1163 467
0 2 39 0 0 8320 0 0 25 64 0 5
1147 395
1197 395
1197 511
1154 511
1154 467
8 4 40 0 0 8320 0 25 25 0 0 5
1136 403
1105 403
1105 477
1136 477
1136 473
3 3 41 0 0 8320 0 25 24 0 0 3
1145 473
1145 511
1095 511
8 4 40 0 0 0 0 25 26 0 0 3
1136 403
1138 403
1138 386
7 3 39 0 0 0 0 25 26 0 0 3
1145 403
1147 403
1147 386
6 2 42 0 0 8320 0 25 26 0 0 3
1154 403
1156 403
1156 386
5 1 19 0 0 0 0 25 26 0 0 3
1163 403
1165 403
1165 386
1 13 43 0 0 8320 0 28 26 0 0 3
1129 292
1111 292
1111 316
2 12 44 0 0 12416 0 28 26 0 0 4
1135 292
1135 297
1120 297
1120 316
3 11 45 0 0 12416 0 28 26 0 0 4
1141 292
1141 301
1129 301
1129 316
4 10 46 0 0 12416 0 28 26 0 0 4
1147 292
1147 303
1138 303
1138 316
5 9 47 0 0 8320 0 28 26 0 0 6
1153 292
1154 292
1154 304
1149 304
1149 316
1147 316
6 8 48 0 0 4224 0 28 26 0 0 3
1159 292
1159 316
1156 316
7 7 49 0 0 4224 0 28 26 0 0 2
1165 292
1165 316
1 2 3 0 0 0 0 27 32 0 0 4
1152 131
1152 150
1151 150
1151 158
1 9 50 0 0 4224 0 32 28 0 0 4
1151 194
1151 212
1150 212
1150 220
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
470 872 618 895
482 882 622 897
20 MODI OMKAR 19EE30018
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
