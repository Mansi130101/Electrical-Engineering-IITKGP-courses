CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 40 10 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
26
9 2-In AND~
219 270 598 0 3 22
0 5 4 6
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U9D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 1798736149
65 0 0 0 4 4 4 0
1 U
8953 0 0
0
0
9 2-In AND~
219 496 619 0 3 22
0 4 5 7
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U9C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
4441 0 0
0
0
8 2-In OR~
219 522 551 0 3 22
0 7 10 11
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U10A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1698072859
65 0 0 0 4 1 5 0
1 U
3618 0 0
0
0
9 2-In AND~
219 553 616 0 3 22
0 9 8 10
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U9B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
6153 0 0
0
0
7 Ground~
168 360 347 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
6 74LS93
109 271 380 0 8 17
0 55 6 8 15 56 57 4 15
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U8
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
6 74LS47
187 237 293 0 14 29
0 2 2 4 15 58 59 22 21 20
19 18 17 16 60
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
2 +V
167 263 75 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V7
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
9 CA 7-Seg~
184 261 187 0 18 19
10 16 17 18 19 20 21 22 61 23
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3549 0 0
0
0
9 CA 7-Seg~
184 516 191 0 18 19
10 25 26 27 28 29 30 31 62 32
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7931 0 0
0
0
2 +V
167 518 79 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
6 74LS47
187 492 297 0 14 29
0 8 5 9 24 63 64 31 30 29
28 27 26 25 65
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U6
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
6 74LS93
109 526 384 0 8 17
0 66 11 12 24 8 5 9 24
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U5
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
6 74LS93
109 764 379 0 8 17
0 12 13 14 33 34 12 13 33
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U4
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
6 74LS47
187 730 292 0 14 29
0 34 12 13 33 67 68 41 40 39
38 37 36 35 69
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
2 +V
167 756 74 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
9 CA 7-Seg~
184 754 186 0 18 19
10 35 36 37 38 39 40 41 70 42
0 0 0 0 2 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3874 0 0
0
0
9 CA 7-Seg~
184 1011 185 0 18 19
10 47 48 49 50 51 52 53 71 54
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6671 0 0
0
0
2 +V
167 1013 73 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
6 74LS47
187 987 291 0 14 29
0 14 46 43 44 72 73 53 52 51
50 49 48 47 74
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
6 74LS93
109 1021 378 0 8 17
0 14 43 45 44 14 46 43 44
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
7 Pulser~
4 923 457 0 10 12
0 75 76 45 77 0 0 5 5 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8778 0 0
0
0
9 Resistor~
219 262 120 0 4 5
0 23 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 517 124 0 4 5
0 32 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 755 119 0 4 5
0 42 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 1012 118 0 4 5
0 54 3 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
76
0 2 4 0 0 4096 0 0 1 5 0 3
334 667
278 667
278 619
0 1 5 0 0 8192 0 0 1 6 0 4
513 668
513 694
260 694
260 619
3 2 6 0 0 4224 0 1 6 0 0 2
269 574
269 410
3 0 7 0 0 8192 0 2 0 0 10 3
495 595
495 597
495 583
0 1 4 0 0 8320 0 0 2 21 0 5
260 338
334 338
334 669
486 669
486 640
2 2 5 0 0 8320 0 12 2 0 0 5
524 334
616 334
616 668
504 668
504 640
0 2 8 0 0 8192 0 0 4 33 0 5
533 343
595 343
595 642
561 642
561 637
0 1 9 0 0 8320 0 0 4 35 0 5
515 340
603 340
603 650
543 650
543 637
2 3 10 0 0 12416 0 3 4 0 0 5
534 567
533 567
533 583
552 583
552 592
1 0 7 0 0 12416 0 3 0 0 0 5
516 567
515 567
515 583
495 583
495 590
2 3 11 0 0 4224 0 13 3 0 0 4
524 414
524 522
525 522
525 521
1 0 2 0 0 4096 0 7 0 0 13 3
278 330
360 330
360 334
2 1 2 0 0 8320 0 7 5 0 0 4
269 330
269 334
360 334
360 341
0 3 12 0 0 8320 0 0 13 16 0 4
791 419
791 467
515 467
515 420
3 0 8 0 0 8320 0 6 0 0 33 5
260 416
260 508
588 508
588 349
533 349
0 1 12 0 0 0 0 0 14 48 0 5
762 338
803 338
803 419
771 419
771 409
0 0 13 0 0 4096 0 0 0 18 18 2
762 333
753 333
2 0 13 0 0 12416 0 14 0 0 49 5
762 409
762 438
829 438
829 333
753 333
0 3 14 0 0 12416 0 0 14 64 0 5
1028 336
1147 336
1147 503
753 503
753 415
4 0 15 0 0 12416 0 6 0 0 22 5
251 416
251 422
226 422
226 338
251 338
3 7 4 0 0 0 0 7 6 0 0 2
260 330
260 346
4 8 15 0 0 0 0 7 6 0 0 2
251 330
251 346
1 13 16 0 0 12416 0 9 7 0 0 4
240 223
240 234
224 234
224 260
2 12 17 0 0 12416 0 9 7 0 0 4
246 223
246 239
233 239
233 260
3 11 18 0 0 4224 0 9 7 0 0 4
252 223
252 244
242 244
242 260
4 10 19 0 0 4224 0 9 7 0 0 4
258 223
258 248
251 248
251 260
5 9 20 0 0 4224 0 9 7 0 0 4
264 223
264 252
260 252
260 260
6 8 21 0 0 4224 0 9 7 0 0 3
270 223
270 260
269 260
7 7 22 0 0 4224 0 9 7 0 0 4
276 223
276 245
278 245
278 260
1 9 23 0 0 8320 0 23 9 0 0 3
262 138
261 138
261 151
1 2 3 0 0 8320 0 8 23 0 0 3
263 84
262 84
262 102
4 0 24 0 0 12416 0 13 0 0 36 5
506 420
506 426
481 426
481 342
506 342
1 5 8 0 0 0 0 12 13 0 0 2
533 334
533 350
2 6 5 0 0 0 0 12 13 0 0 2
524 334
524 350
3 7 9 0 0 0 0 12 13 0 0 2
515 334
515 350
4 8 24 0 0 0 0 12 13 0 0 2
506 334
506 350
1 13 25 0 0 12416 0 10 12 0 0 4
495 227
495 238
479 238
479 264
2 12 26 0 0 12416 0 10 12 0 0 4
501 227
501 243
488 243
488 264
3 11 27 0 0 4224 0 10 12 0 0 4
507 227
507 248
497 248
497 264
4 10 28 0 0 4224 0 10 12 0 0 4
513 227
513 252
506 252
506 264
5 9 29 0 0 4224 0 10 12 0 0 4
519 227
519 256
515 256
515 264
6 8 30 0 0 4224 0 10 12 0 0 3
525 227
525 264
524 264
7 7 31 0 0 4224 0 10 12 0 0 4
531 227
531 249
533 249
533 264
1 9 32 0 0 8320 0 24 10 0 0 3
517 142
516 142
516 155
1 2 3 0 0 0 0 11 24 0 0 3
518 88
517 88
517 106
4 0 33 0 0 12416 0 14 0 0 50 5
744 415
744 421
719 421
719 337
744 337
1 5 34 0 0 4224 0 15 14 0 0 2
771 329
771 345
2 6 12 0 0 0 0 15 14 0 0 2
762 329
762 345
3 7 13 0 0 0 0 15 14 0 0 2
753 329
753 345
4 8 33 0 0 0 0 15 14 0 0 2
744 329
744 345
1 13 35 0 0 12416 0 17 15 0 0 4
733 222
733 233
717 233
717 259
2 12 36 0 0 12416 0 17 15 0 0 4
739 222
739 238
726 238
726 259
3 11 37 0 0 4224 0 17 15 0 0 4
745 222
745 243
735 243
735 259
4 10 38 0 0 4224 0 17 15 0 0 4
751 222
751 247
744 247
744 259
5 9 39 0 0 4224 0 17 15 0 0 4
757 222
757 251
753 251
753 259
6 8 40 0 0 4224 0 17 15 0 0 3
763 222
763 259
762 259
7 7 41 0 0 4224 0 17 15 0 0 4
769 222
769 244
771 244
771 259
1 9 42 0 0 8320 0 25 17 0 0 3
755 137
754 137
754 150
1 2 3 0 0 0 0 16 25 0 0 3
756 83
755 83
755 101
1 5 14 0 0 0 0 21 21 0 0 5
1028 408
1028 430
1073 430
1073 344
1028 344
3 2 43 0 0 8320 0 20 21 0 0 5
1010 328
1095 328
1095 446
1019 446
1019 408
4 0 44 0 0 12416 0 21 0 0 67 5
1001 414
1001 420
976 420
976 336
1001 336
3 3 45 0 0 4224 0 22 21 0 0 3
947 448
1010 448
1010 414
1 5 14 0 0 0 0 20 21 0 0 2
1028 328
1028 344
2 6 46 0 0 4224 0 20 21 0 0 2
1019 328
1019 344
3 7 43 0 0 0 0 20 21 0 0 2
1010 328
1010 344
4 8 44 0 0 0 0 20 21 0 0 2
1001 328
1001 344
1 13 47 0 0 12416 0 18 20 0 0 4
990 221
990 232
974 232
974 258
2 12 48 0 0 12416 0 18 20 0 0 4
996 221
996 237
983 237
983 258
3 11 49 0 0 4224 0 18 20 0 0 4
1002 221
1002 242
992 242
992 258
4 10 50 0 0 4224 0 18 20 0 0 4
1008 221
1008 246
1001 246
1001 258
5 9 51 0 0 4224 0 18 20 0 0 4
1014 221
1014 250
1010 250
1010 258
6 8 52 0 0 4224 0 18 20 0 0 3
1020 221
1020 258
1019 258
7 7 53 0 0 4224 0 18 20 0 0 4
1026 221
1026 243
1028 243
1028 258
1 9 54 0 0 8320 0 26 18 0 0 3
1012 136
1011 136
1011 149
1 2 3 0 0 0 0 19 26 0 0 3
1013 82
1012 82
1012 100
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2361676 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
4720856 8419392 100 100 0 0
77 66 1487 276
0 447 1536 823
1487 66
77 66
1487 66
1487 276
0 0
4.53041e-315 0 4.53041e-315 0 4.53041e-315 4.53041e-315
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
