CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 1 80 9
0 70 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1280 680
177209362 0
0
6 Title:
5 Name:
0
0
0
22
9 2-In AND~
219 113 466 0 3 22
0 3 4 5
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U7C
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 5 0
1 U
8953 0 0
0
0
8 2-In OR~
219 71 504 0 3 22
0 5 6 7
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U8A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2010083361
65 0 0 0 4 1 6 0
1 U
4441 0 0
0
0
9 2-In AND~
219 43 344 0 3 22
0 3 9 8
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U7B
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
3618 0 0
0
0
9 2-In AND~
219 67 299 0 3 22
0 10 9 6
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U7A
4 13 25 21
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
6153 0 0
0
0
8 3-In OR~
219 23 457 0 4 22
0 6 8 4 11
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U6C
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 4 0
1 U
5394 0 0
0
0
9 2-In AND~
219 107 299 0 3 22
0 3 4 13
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U4D
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
7734 0 0
0
0
9 2-In AND~
219 146 299 0 3 22
0 10 3 14
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U4C
5 18 26 26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
9914 0 0
0
0
8 3-In OR~
219 178 459 0 4 22
0 6 14 13 12
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U6B
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 4 0
1 U
3747 0 0
0
0
8 3-In OR~
219 224 424 0 4 22
0 16 17 18 15
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U6A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3549 0 0
0
0
9 3-In AND~
219 177 346 0 4 22
0 19 10 3 18
0
0 0 608 270
6 74LS11
-21 -28 21 -20
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
7931 0 0
0
0
9 2-In AND~
219 230 349 0 3 22
0 20 21 17
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9325 0 0
0
0
9 2-In AND~
219 285 347 0 3 22
0 9 20 16
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2093969452
65 0 0 0 4 1 2 0
1 U
8903 0 0
0
0
9 Inverter~
13 303 240 0 2 22
0 19 9
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U3C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
3834 0 0
0
0
9 Inverter~
13 256 239 0 2 22
0 10 20
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U3B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
3363 0 0
0
0
9 Inverter~
13 202 240 0 2 22
0 3 21
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
7668 0 0
0
0
7 Pulser~
4 69 98 0 10 12
0 33 34 35 22 0 0 5 5 6
7
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
6 74LS90
107 182 145 0 10 21
0 2 36 37 2 22 3 4 19 10
3
0
0 0 13024 270
6 74LS90
-21 -51 21 -43
2 U2
40 -4 54 4
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
7 Ground~
168 175 91 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
9 CA 7-Seg~
184 68 640 0 18 19
10 25 26 27 28 30 29 31 38 24
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-62 -24 -27 -16
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3789 0 0
0
0
2 +V
167 68 560 0 1 3
0 23
0
0 0 54240 0
2 5V
-29 13 -15 21
2 V1
-27 2 -13 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4871 0 0
0
0
6 74LS47
187 186 637 0 14 29
0 11 7 12 15 39 40 31 29 30
28 27 26 25 41
0
0 0 13024 782
6 74LS47
-21 -60 21 -52
2 U1
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
9 Resistor~
219 68 587 0 4 5
0 24 23 0 1
0
0 0 864 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
48
1 1 3 0 0 4096 0 1 3 0 0 4
120 444
120 347
50 347
50 322
2 0 4 0 0 12288 0 1 0 0 13 4
102 444
97 444
97 396
17 396
3 1 5 0 0 8320 0 1 2 0 0 4
111 489
111 487
83 487
83 488
2 0 6 0 0 4096 0 2 0 0 9 2
65 488
65 420
3 2 7 0 0 8320 0 2 21 0 0 4
74 534
74 533
160 533
160 604
1 0 3 0 0 0 0 3 0 0 17 4
50 322
45 322
45 258
114 258
3 2 8 0 0 8320 0 3 5 0 0 3
41 367
26 367
26 442
2 0 9 0 0 4096 0 3 0 0 11 3
32 322
32 266
56 266
1 0 6 0 0 0 0 5 0 0 12 3
35 441
35 420
65 420
1 0 10 0 0 8192 0 4 0 0 21 3
74 277
74 248
158 248
2 0 9 0 0 8320 0 4 0 0 31 3
56 277
56 266
306 266
3 1 6 0 0 8320 0 4 8 0 0 4
65 322
65 420
190 420
190 443
3 0 4 0 0 4224 0 5 0 0 16 3
17 441
17 232
96 232
4 1 11 0 0 8320 0 5 21 0 0 4
26 487
26 540
151 540
151 604
4 3 12 0 0 8320 0 8 21 0 0 3
181 489
169 489
169 604
2 7 4 0 0 0 0 6 17 0 0 4
96 277
96 184
202 184
202 178
1 0 3 0 0 0 0 6 0 0 20 3
114 277
114 257
135 257
3 3 13 0 0 4224 0 6 8 0 0 4
105 322
105 437
172 437
172 443
3 2 14 0 0 4224 0 7 8 0 0 4
144 322
144 428
181 428
181 444
2 0 3 0 0 0 0 7 0 0 35 3
135 277
135 200
148 200
1 0 10 0 0 0 0 7 0 0 34 4
153 277
158 277
158 199
166 199
4 4 15 0 0 4224 0 9 21 0 0 4
227 454
227 596
178 596
178 604
1 3 16 0 0 8320 0 9 12 0 0 4
236 408
236 378
283 378
283 370
2 3 17 0 0 4224 0 9 11 0 0 4
227 409
227 380
228 380
228 372
3 4 18 0 0 8320 0 9 10 0 0 4
218 408
218 376
175 376
175 369
1 0 19 0 0 4224 0 10 0 0 33 2
184 324
184 189
2 0 10 0 0 4224 0 10 0 0 34 2
175 324
175 201
3 0 3 0 0 4224 0 10 0 0 35 2
166 324
166 214
2 1 20 0 0 8320 0 14 11 0 0 5
259 257
255 257
255 319
237 319
237 327
2 2 21 0 0 4224 0 15 11 0 0 4
205 258
205 319
219 319
219 327
2 1 9 0 0 0 0 13 12 0 0 4
306 258
306 317
292 317
292 325
2 2 20 0 0 0 0 14 12 0 0 5
259 257
262 257
262 317
274 317
274 325
8 1 19 0 0 0 0 17 13 0 0 4
184 178
184 189
306 189
306 222
9 1 10 0 0 0 0 17 14 0 0 4
166 178
166 201
259 201
259 221
10 1 3 0 0 0 0 17 15 0 0 4
148 178
148 214
205 214
205 222
1 0 2 0 0 0 0 18 0 0 37 2
175 99
175 99
4 1 2 0 0 8320 0 17 17 0 0 4
175 114
175 99
202 99
202 114
6 10 3 0 0 0 0 17 17 0 0 6
148 108
148 103
134 103
134 177
148 177
148 178
4 5 22 0 0 4224 0 16 17 0 0 3
99 98
157 98
157 108
1 2 23 0 0 0 0 20 22 0 0 2
68 569
68 569
1 9 24 0 0 4224 0 22 19 0 0 2
68 605
68 604
1 13 25 0 0 8320 0 19 21 0 0 4
47 676
47 685
205 685
205 674
12 2 26 0 0 8320 0 21 19 0 0 4
196 674
196 684
53 684
53 676
11 3 27 0 0 8320 0 21 19 0 0 4
187 674
187 684
59 684
59 676
10 4 28 0 0 8320 0 21 19 0 0 4
178 674
178 684
65 684
65 676
8 6 29 0 0 8320 0 21 19 0 0 4
160 674
160 684
77 684
77 676
9 5 30 0 0 8320 0 21 19 0 0 4
169 674
169 684
71 684
71 676
7 7 31 0 0 8320 0 21 19 0 0 4
151 674
151 684
83 684
83 676
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
512 118 616 182
522 126 618 174
23 MANSI UNIYAL
19EE10039
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 152
481 187 699 324
494 197 704 302
152 roll number dsiplay using 
counter and logic gates:

E will be displayed by symbol 
display of 14
and last letter will be blank 
and then reset
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
5703132 1079360 100 100 0 0
0 0 0 0
267 81 428 151
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2622868 8419392 100 100 0 0
77 66 1007 216
267 385 1308 689
1007 66
77 66
1007 66
1007 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
