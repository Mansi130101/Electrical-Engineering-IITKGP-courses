CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 294 69 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-38 -17 -24 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3226 0 0
2
44497.7 0
0
7 Pulser~
4 142 50 0 10 12
0 47 48 3 49 0 0 5 5 1
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6966 0 0
2
44497.7 0
0
2 +V
167 350 309 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9796 0 0
2
44497.7 0
0
2 +V
167 692 409 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5952 0 0
2
5.90006e-315 0
0
9 CA 7-Seg~
184 762 538 0 18 19
10 14 13 12 11 10 9 8 50 6
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3649 0 0
2
5.90006e-315 0
0
9 CA 7-Seg~
184 615 538 0 18 19
10 21 20 19 18 17 16 15 51 7
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3716 0 0
2
5.90006e-315 0
0
6 74LS47
187 401 537 0 14 29
0 25 23 24 22 52 53 8 9 10
11 12 13 14 54
0
0 0 4848 270
6 74LS47
-21 -60 21 -52
2 U6
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4797 0 0
2
5.90006e-315 0
0
6 74LS47
187 246 535 0 14 29
0 29 28 27 26 55 56 15 16 17
18 19 20 21 57
0
0 0 4848 270
6 74LS47
-21 -60 21 -52
2 U5
60 -5 74 3
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4681 0 0
2
5.90006e-315 0
0
6 74LS83
105 430 327 0 14 29
0 38 37 36 35 42 41 40 39 4
25 23 24 22 30
0
0 0 4848 270
5 74F83
-18 -60 17 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9730 0 0
2
5.90006e-315 0
0
6 74LS83
105 276 329 0 14 29
0 34 33 32 31 46 45 44 43 30
29 28 27 26 58
0
0 0 4848 270
5 74F83
-18 -60 17 -52
2 U3
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
9874 0 0
2
5.90006e-315 0
0
7 74LS273
150 468 150 0 18 37
0 2 3 39 40 41 42 43 44 45
46 35 36 37 38 31 32 33 34
0
0 0 4848 692
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
364 0 0
2
5.90006e-315 0
0
7 74LS273
150 252 150 0 18 37
0 2 3 22 24 23 25 26 27 28
29 39 40 41 42 43 44 45 46
0
0 0 4848 692
7 74LS273
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3656 0 0
2
5.90006e-315 0
0
9 Resistor~
219 762 467 0 4 5
0 6 5 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3131 0 0
2
5.90006e-315 0
0
9 Resistor~
219 615 467 0 4 5
0 7 5 0 1
0
0 0 880 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6772 0 0
2
5.90006e-315 0
0
64
1 1 2 0 0 8320 0 1 11 0 0 4
294 81
294 90
430 90
430 190
1 1 2 0 0 16 0 1 12 0 0 6
294 81
340 81
340 210
206 210
206 190
214 190
3 2 3 0 0 4224 0 2 11 0 0 4
166 41
422 41
422 181
436 181
3 2 3 0 0 0 0 2 12 0 0 4
166 41
209 41
209 181
220 181
1 9 4 0 0 12416 0 3 9 0 0 6
350 318
350 317
373 317
373 292
387 292
387 297
1 2 5 0 0 4096 0 4 13 0 0 3
692 418
762 418
762 449
2 1 5 0 0 8320 0 14 4 0 0 3
615 449
615 418
692 418
9 1 6 0 0 4224 0 5 13 0 0 2
762 502
762 485
9 1 7 0 0 4224 0 6 14 0 0 2
615 502
615 485
7 7 8 0 0 8320 0 7 5 0 0 4
442 574
442 772
777 772
777 574
6 8 9 0 0 8320 0 5 7 0 0 4
771 574
771 759
433 759
433 574
9 5 10 0 0 8320 0 7 5 0 0 4
424 574
424 747
765 747
765 574
4 10 11 0 0 8320 0 5 7 0 0 4
759 574
759 736
415 736
415 574
11 3 12 0 0 8320 0 7 5 0 0 4
406 574
406 725
753 725
753 574
2 12 13 0 0 8320 0 5 7 0 0 4
747 574
747 708
397 708
397 574
13 1 14 0 0 8320 0 7 5 0 0 4
388 574
388 716
741 716
741 574
7 7 15 0 0 8320 0 8 6 0 0 4
287 572
287 661
630 661
630 574
6 8 16 0 0 8320 0 6 8 0 0 4
624 574
624 648
278 648
278 572
9 5 17 0 0 8320 0 8 6 0 0 4
269 572
269 636
618 636
618 574
4 10 18 0 0 8320 0 6 8 0 0 4
612 574
612 625
260 625
260 572
11 3 19 0 0 8320 0 8 6 0 0 4
251 572
251 614
606 614
606 574
2 12 20 0 0 8320 0 6 8 0 0 4
600 574
600 597
242 597
242 572
13 1 21 0 0 8320 0 8 6 0 0 4
233 572
233 605
594 605
594 574
3 0 22 0 0 8320 0 12 0 0 32 4
220 172
175 172
175 449
414 449
0 5 23 0 0 8320 0 0 12 34 0 4
432 467
150 467
150 154
220 154
4 0 24 0 0 8320 0 12 0 0 33 4
220 163
162 163
162 458
423 458
6 0 25 0 0 8320 0 12 0 0 35 4
220 145
139 145
139 478
441 478
7 0 26 0 0 8320 0 12 0 0 36 4
220 136
127 136
127 396
260 396
0 8 27 0 0 8320 0 0 12 37 0 4
269 407
116 407
116 127
220 127
9 0 28 0 0 8320 0 12 0 0 38 4
220 118
104 118
104 416
278 416
10 0 29 0 0 8320 0 12 0 0 39 4
220 109
91 109
91 424
287 424
13 4 22 0 0 0 0 9 7 0 0 4
414 361
414 449
415 449
415 504
3 12 24 0 0 0 0 7 9 0 0 4
424 504
424 458
423 458
423 361
11 2 23 0 0 0 0 9 7 0 0 4
432 361
432 467
433 467
433 504
10 1 25 0 0 0 0 9 7 0 0 4
441 361
441 478
442 478
442 504
13 4 26 0 0 0 0 10 8 0 0 2
260 363
260 502
3 12 27 0 0 0 0 8 10 0 0 2
269 502
269 363
11 2 28 0 0 0 0 10 8 0 0 2
278 363
278 502
10 1 29 0 0 0 0 10 8 0 0 2
287 363
287 502
9 14 30 0 0 16512 0 10 9 0 0 6
233 299
233 286
194 286
194 382
387 382
387 361
15 4 31 0 0 12416 0 11 10 0 0 5
500 136
566 136
566 262
287 262
287 299
3 16 32 0 0 8320 0 10 11 0 0 5
296 299
296 270
576 270
576 127
500 127
17 2 33 0 0 12416 0 11 10 0 0 5
500 118
584 118
584 278
305 278
305 299
1 18 34 0 0 8320 0 10 11 0 0 5
314 299
314 286
594 286
594 109
500 109
11 4 35 0 0 12416 0 11 9 0 0 5
500 172
514 172
514 229
441 229
441 297
3 12 36 0 0 12416 0 9 11 0 0 5
450 297
450 237
523 237
523 163
500 163
13 2 37 0 0 8320 0 11 9 0 0 5
500 154
530 154
530 244
459 244
459 297
1 14 38 0 0 12416 0 9 11 0 0 5
468 297
468 255
540 255
540 145
500 145
0 8 39 0 0 4096 0 0 9 57 0 4
359 172
359 250
405 250
405 297
7 0 40 0 0 12288 0 9 0 0 58 4
414 297
414 244
367 244
367 163
0 6 41 0 0 4096 0 0 9 59 0 4
375 154
375 235
423 235
423 297
5 0 42 0 0 12288 0 9 0 0 60 4
432 297
432 227
385 227
385 145
0 8 43 0 0 4096 0 0 10 61 0 4
294 136
294 221
251 221
251 299
7 0 44 0 0 12288 0 10 0 0 62 4
260 299
260 230
302 230
302 127
6 0 45 0 0 12288 0 10 0 0 63 4
269 299
269 237
311 237
311 118
5 0 46 0 0 12288 0 10 0 0 64 4
278 299
278 245
323 245
323 109
11 3 39 0 0 4224 0 12 11 0 0 2
284 172
436 172
4 12 40 0 0 4224 0 11 12 0 0 2
436 163
284 163
13 5 41 0 0 4224 0 12 11 0 0 2
284 154
436 154
6 14 42 0 0 4224 0 11 12 0 0 2
436 145
284 145
15 7 43 0 0 4224 0 12 11 0 0 2
284 136
436 136
8 16 44 0 0 4224 0 11 12 0 0 2
436 127
284 127
17 9 45 0 0 4224 0 12 11 0 0 2
284 118
436 118
18 10 46 0 0 4224 0 12 11 0 0 2
284 109
436 109
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
